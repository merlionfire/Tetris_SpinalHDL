// Generator : SpinalHDL dev    git head : f518b561b4631c190dbd783ec02e46e2c7fbf8ff
// Component : top
// Git hash  : f549e498c0dad121e3d5ad08cc969073c9d4a436

`timescale 1ns/1ps

module top (
  output              io_vga_vSync,
  output              io_vga_hSync,
  output              io_vga_colorEn,
  output     [3:0]    io_vga_color_r,
  output     [3:0]    io_vga_color_g,
  output     [3:0]    io_vga_color_b,
  input               io_patgen_sel,
  input               clk,
  input               reset
);

  wire                patgen_1_io_sel;
  wire                objects_io_inside;
  wire       [3:0]    objects_io_color_r;
  wire       [3:0]    objects_io_color_g;
  wire       [3:0]    objects_io_color_b;
  wire       [3:0]    patgen_1_io_color_r;
  wire       [3:0]    patgen_1_io_color_g;
  wire       [3:0]    patgen_1_io_color_b;
  wire                ctrl_io_frameStart;
  wire                ctrl_io_pixels_ready;
  wire                ctrl_io_vga_vSync;
  wire                ctrl_io_vga_hSync;
  wire                ctrl_io_vga_colorEn;
  wire       [3:0]    ctrl_io_vga_color_r;
  wire       [3:0]    ctrl_io_vga_color_g;
  wire       [3:0]    ctrl_io_vga_color_b;
  wire                ctrl_io_error;
  reg        [9:0]    x_addr;
  reg        [9:0]    y_addr;
  reg                 toplevel_ctrl_io_vga_colorEn_regNext;
  wire                when_top_l36;
  reg                 io_patgen_sel_regNext;

  layout objects (
    .io_x       (x_addr[9:0]            ), //i
    .io_y       (y_addr[9:0]            ), //i
    .io_inside  (objects_io_inside      ), //o
    .io_color_r (objects_io_color_r[3:0]), //o
    .io_color_g (objects_io_color_g[3:0]), //o
    .io_color_b (objects_io_color_b[3:0]), //o
    .clk        (clk                    ), //i
    .reset      (reset                  )  //i
  );
  patgen patgen_1 (
    .io_color_en (ctrl_io_vga_colorEn     ), //i
    .io_x        (x_addr[9:0]             ), //i
    .io_y        (y_addr[9:0]             ), //i
    .io_sel      (patgen_1_io_sel         ), //i
    .io_color_r  (patgen_1_io_color_r[3:0]), //o
    .io_color_g  (patgen_1_io_color_g[3:0]), //o
    .io_color_b  (patgen_1_io_color_b[3:0]), //o
    .clk         (clk                     ), //i
    .reset       (reset                   )  //i
  );
  VgaCtrl ctrl (
    .io_softReset            (1'b0                    ), //i
    .io_timings_h_syncStart  (11'h087                 ), //i
    .io_timings_h_syncEnd    (11'h52f                 ), //i
    .io_timings_h_colorStart (11'h117                 ), //i
    .io_timings_h_colorEnd   (11'h517                 ), //i
    .io_timings_h_polarity   (1'b0                    ), //i
    .io_timings_v_syncStart  (11'h005                 ), //i
    .io_timings_v_syncEnd    (11'h325                 ), //i
    .io_timings_v_colorStart (11'h022                 ), //i
    .io_timings_v_colorEnd   (11'h322                 ), //i
    .io_timings_v_polarity   (1'b0                    ), //i
    .io_frameStart           (ctrl_io_frameStart      ), //o
    .io_pixels_valid         (1'b1                    ), //i
    .io_pixels_ready         (ctrl_io_pixels_ready    ), //o
    .io_pixels_payload_r     (patgen_1_io_color_r[3:0]), //i
    .io_pixels_payload_g     (patgen_1_io_color_g[3:0]), //i
    .io_pixels_payload_b     (patgen_1_io_color_b[3:0]), //i
    .io_vga_vSync            (ctrl_io_vga_vSync       ), //o
    .io_vga_hSync            (ctrl_io_vga_hSync       ), //o
    .io_vga_colorEn          (ctrl_io_vga_colorEn     ), //o
    .io_vga_color_r          (ctrl_io_vga_color_r[3:0]), //o
    .io_vga_color_g          (ctrl_io_vga_color_g[3:0]), //o
    .io_vga_color_b          (ctrl_io_vga_color_b[3:0]), //o
    .io_error                (ctrl_io_error           ), //o
    .clk                     (clk                     ), //i
    .reset                   (reset                   )  //i
  );
  assign when_top_l36 = ((! ctrl_io_vga_colorEn) && toplevel_ctrl_io_vga_colorEn_regNext);
  assign patgen_1_io_sel = (io_patgen_sel && (! io_patgen_sel_regNext));
  assign io_vga_vSync = ctrl_io_vga_vSync;
  assign io_vga_hSync = ctrl_io_vga_hSync;
  assign io_vga_colorEn = ctrl_io_vga_colorEn;
  assign io_vga_color_r = ctrl_io_vga_color_r;
  assign io_vga_color_g = ctrl_io_vga_color_g;
  assign io_vga_color_b = ctrl_io_vga_color_b;
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      x_addr <= 10'h0;
      y_addr <= 10'h0;
      io_patgen_sel_regNext <= 1'b0;
    end else begin
      if(ctrl_io_vga_colorEn) begin
        x_addr <= (x_addr + 10'h001);
      end else begin
        x_addr <= 10'h0;
      end
      if(ctrl_io_frameStart) begin
        y_addr <= 10'h0;
      end else begin
        if(when_top_l36) begin
          y_addr <= (y_addr + 10'h001);
        end
      end
      io_patgen_sel_regNext <= io_patgen_sel;
    end
  end

  always @(posedge clk) begin
    toplevel_ctrl_io_vga_colorEn_regNext <= ctrl_io_vga_colorEn;
  end


endmodule

module VgaCtrl (
  input               io_softReset,
  input      [10:0]   io_timings_h_syncStart,
  input      [10:0]   io_timings_h_syncEnd,
  input      [10:0]   io_timings_h_colorStart,
  input      [10:0]   io_timings_h_colorEnd,
  input               io_timings_h_polarity,
  input      [10:0]   io_timings_v_syncStart,
  input      [10:0]   io_timings_v_syncEnd,
  input      [10:0]   io_timings_v_colorStart,
  input      [10:0]   io_timings_v_colorEnd,
  input               io_timings_v_polarity,
  output              io_frameStart,
  input               io_pixels_valid,
  output              io_pixels_ready,
  input      [3:0]    io_pixels_payload_r,
  input      [3:0]    io_pixels_payload_g,
  input      [3:0]    io_pixels_payload_b,
  output              io_vga_vSync,
  output              io_vga_hSync,
  output              io_vga_colorEn,
  output     [3:0]    io_vga_color_r,
  output     [3:0]    io_vga_color_g,
  output     [3:0]    io_vga_color_b,
  output              io_error,
  input               clk,
  input               reset
);

  wire                when_VgaCtrl_l183;
  reg        [10:0]   h_counter;
  wire                h_syncStart;
  wire                h_syncEnd;
  wire                h_colorStart;
  wire                h_colorEnd;
  reg                 h_sync;
  reg                 h_colorEn;
  reg        [10:0]   v_counter;
  wire                v_syncStart;
  wire                v_syncEnd;
  wire                v_colorStart;
  wire                v_colorEnd;
  reg                 v_sync;
  reg                 v_colorEn;
  wire                colorEn;

  assign when_VgaCtrl_l183 = 1'b1;
  assign h_syncStart = (h_counter == io_timings_h_syncStart);
  assign h_syncEnd = (h_counter == io_timings_h_syncEnd);
  assign h_colorStart = (h_counter == io_timings_h_colorStart);
  assign h_colorEnd = (h_counter == io_timings_h_colorEnd);
  assign v_syncStart = (v_counter == io_timings_v_syncStart);
  assign v_syncEnd = (v_counter == io_timings_v_syncEnd);
  assign v_colorStart = (v_counter == io_timings_v_colorStart);
  assign v_colorEnd = (v_counter == io_timings_v_colorEnd);
  assign colorEn = (h_colorEn && v_colorEn);
  assign io_pixels_ready = colorEn;
  assign io_error = (colorEn && (! io_pixels_valid));
  assign io_frameStart = (v_syncStart && h_syncStart);
  assign io_vga_hSync = (h_sync ^ io_timings_h_polarity);
  assign io_vga_vSync = (v_sync ^ io_timings_v_polarity);
  assign io_vga_colorEn = colorEn;
  assign io_vga_color_r = io_pixels_payload_r;
  assign io_vga_color_g = io_pixels_payload_g;
  assign io_vga_color_b = io_pixels_payload_b;
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      h_counter <= 11'h0;
      h_sync <= 1'b0;
      h_colorEn <= 1'b0;
      v_counter <= 11'h0;
      v_sync <= 1'b0;
      v_colorEn <= 1'b0;
    end else begin
      if(when_VgaCtrl_l183) begin
        h_counter <= (h_counter + 11'h001);
        if(h_syncEnd) begin
          h_counter <= 11'h0;
        end
      end
      if(h_syncStart) begin
        h_sync <= 1'b1;
      end
      if(h_syncEnd) begin
        h_sync <= 1'b0;
      end
      if(h_colorStart) begin
        h_colorEn <= 1'b1;
      end
      if(h_colorEnd) begin
        h_colorEn <= 1'b0;
      end
      if(io_softReset) begin
        h_counter <= 11'h0;
        h_sync <= 1'b0;
        h_colorEn <= 1'b0;
      end
      if(h_syncEnd) begin
        v_counter <= (v_counter + 11'h001);
        if(v_syncEnd) begin
          v_counter <= 11'h0;
        end
      end
      if(v_syncStart) begin
        v_sync <= 1'b1;
      end
      if(v_syncEnd) begin
        v_sync <= 1'b0;
      end
      if(v_colorStart) begin
        v_colorEn <= 1'b1;
      end
      if(v_colorEnd) begin
        v_colorEn <= 1'b0;
      end
      if(io_softReset) begin
        v_counter <= 11'h0;
        v_sync <= 1'b0;
        v_colorEn <= 1'b0;
      end
    end
  end


endmodule

module patgen (
  input               io_color_en,
  input      [9:0]    io_x,
  input      [9:0]    io_y,
  input               io_sel,
  output     [3:0]    io_color_r,
  output     [3:0]    io_color_g,
  output     [3:0]    io_color_b,
  input               clk,
  input               reset
);

  wire       [1:0]    _zz_sel_id_valueNext;
  wire       [0:0]    _zz_sel_id_valueNext_1;
  wire       [3:0]    _zz_color_bar_idx;
  wire       [5:0]    _zz_color_palette_idx;
  wire       [5:0]    _zz_color_palette_idx_1;
  wire       [5:0]    _zz_color_palette_idx_2;
  wire       [5:0]    _zz_color_palette_idx_3;
  reg                 sel_id_willIncrement;
  wire                sel_id_willClear;
  reg        [1:0]    sel_id_valueNext;
  reg        [1:0]    sel_id_value;
  wire                sel_id_willOverflowIfInc;
  wire                sel_id_willOverflow;
  wire       [3:0]    color_blank_r;
  wire       [3:0]    color_blank_g;
  wire       [3:0]    color_blank_b;
  reg        [3:0]    color_bar_color_r;
  reg        [3:0]    color_bar_color_g;
  reg        [3:0]    color_bar_color_b;
  wire       [4:0]    color_bar_idx;
  reg        [3:0]    color_palette_color_r;
  wire       [3:0]    color_palette_color_g;
  wire       [3:0]    color_palette_color_b;
  wire       [11:0]   color_palette_idx;
  wire       [3:0]    color_palette_color_vec_0;
  wire       [3:0]    color_palette_color_vec_1;
  wire       [3:0]    color_palette_color_vec_2;
  wire                when_patgen_l87;
  reg        [3:0]    _zz_io_color_r;
  reg        [3:0]    _zz_io_color_g;
  reg        [3:0]    _zz_io_color_b;

  assign _zz_sel_id_valueNext_1 = sel_id_willIncrement;
  assign _zz_sel_id_valueNext = {1'd0, _zz_sel_id_valueNext_1};
  assign _zz_color_bar_idx = io_x[9 : 6];
  assign _zz_color_palette_idx_1 = io_y[9 : 4];
  assign _zz_color_palette_idx = _zz_color_palette_idx_1;
  assign _zz_color_palette_idx_3 = io_x[9 : 4];
  assign _zz_color_palette_idx_2 = _zz_color_palette_idx_3;
  always @(*) begin
    sel_id_willIncrement = 1'b0;
    if(io_sel) begin
      sel_id_willIncrement = 1'b1;
    end
  end

  assign sel_id_willClear = 1'b0;
  assign sel_id_willOverflowIfInc = (sel_id_value == 2'b10);
  assign sel_id_willOverflow = (sel_id_willOverflowIfInc && sel_id_willIncrement);
  always @(*) begin
    if(sel_id_willOverflow) begin
      sel_id_valueNext = 2'b00;
    end else begin
      sel_id_valueNext = (sel_id_value + _zz_sel_id_valueNext);
    end
    if(sel_id_willClear) begin
      sel_id_valueNext = 2'b00;
    end
  end

  assign color_blank_r = 4'b0000;
  assign color_blank_g = 4'b0000;
  assign color_blank_b = 4'b0000;
  assign color_bar_idx = {1'd0, _zz_color_bar_idx};
  always @(*) begin
    case(color_bar_idx)
      5'h0 : begin
        color_bar_color_b = 4'b0000;
      end
      5'h01 : begin
        color_bar_color_b = 4'b0111;
      end
      5'h02 : begin
        color_bar_color_b = 4'b1111;
      end
      5'h03 : begin
        color_bar_color_b = 4'b0000;
      end
      5'h04 : begin
        color_bar_color_b = 4'b1111;
      end
      5'h05 : begin
        color_bar_color_b = 4'b1111;
      end
      5'h06 : begin
        color_bar_color_b = 4'b0000;
      end
      5'h07 : begin
        color_bar_color_b = 4'b0111;
      end
      5'h08 : begin
        color_bar_color_b = 4'b1111;
      end
      5'h09 : begin
        color_bar_color_b = 4'b0000;
      end
      5'h0a : begin
        color_bar_color_b = 4'b1111;
      end
      5'h0b : begin
        color_bar_color_b = 4'b1111;
      end
      5'h0c : begin
        color_bar_color_b = 4'b0000;
      end
      5'h0d : begin
        color_bar_color_b = 4'b0111;
      end
      5'h0e : begin
        color_bar_color_b = 4'b1111;
      end
      5'h0f : begin
        color_bar_color_b = 4'b0000;
      end
      5'h10 : begin
        color_bar_color_b = 4'b1111;
      end
      5'h11 : begin
        color_bar_color_b = 4'b1111;
      end
      5'h12 : begin
        color_bar_color_b = 4'b0000;
      end
      5'h13 : begin
        color_bar_color_b = 4'b0101;
      end
      default : begin
        color_bar_color_b = 4'b0000;
      end
    endcase
  end

  always @(*) begin
    case(color_bar_idx)
      5'h0 : begin
        color_bar_color_g = 4'b0000;
      end
      5'h01 : begin
        color_bar_color_g = 4'b0000;
      end
      5'h02 : begin
        color_bar_color_g = 4'b0000;
      end
      5'h03 : begin
        color_bar_color_g = 4'b0111;
      end
      5'h04 : begin
        color_bar_color_g = 4'b0111;
      end
      5'h05 : begin
        color_bar_color_g = 4'b1111;
      end
      5'h06 : begin
        color_bar_color_g = 4'b0000;
      end
      5'h07 : begin
        color_bar_color_g = 4'b0000;
      end
      5'h08 : begin
        color_bar_color_g = 4'b0000;
      end
      5'h09 : begin
        color_bar_color_g = 4'b0111;
      end
      5'h0a : begin
        color_bar_color_g = 4'b0111;
      end
      5'h0b : begin
        color_bar_color_g = 4'b1111;
      end
      5'h0c : begin
        color_bar_color_g = 4'b0000;
      end
      5'h0d : begin
        color_bar_color_g = 4'b0000;
      end
      5'h0e : begin
        color_bar_color_g = 4'b0000;
      end
      5'h0f : begin
        color_bar_color_g = 4'b0111;
      end
      5'h10 : begin
        color_bar_color_g = 4'b0111;
      end
      5'h11 : begin
        color_bar_color_g = 4'b1111;
      end
      5'h12 : begin
        color_bar_color_g = 4'b0101;
      end
      5'h13 : begin
        color_bar_color_g = 4'b0000;
      end
      default : begin
        color_bar_color_g = 4'b0000;
      end
    endcase
  end

  always @(*) begin
    case(color_bar_idx)
      5'h0 : begin
        color_bar_color_r = 4'b1111;
      end
      5'h01 : begin
        color_bar_color_r = 4'b0000;
      end
      5'h02 : begin
        color_bar_color_r = 4'b0000;
      end
      5'h03 : begin
        color_bar_color_r = 4'b0000;
      end
      5'h04 : begin
        color_bar_color_r = 4'b0000;
      end
      5'h05 : begin
        color_bar_color_r = 4'b0000;
      end
      5'h06 : begin
        color_bar_color_r = 4'b0111;
      end
      5'h07 : begin
        color_bar_color_r = 4'b0111;
      end
      5'h08 : begin
        color_bar_color_r = 4'b0111;
      end
      5'h09 : begin
        color_bar_color_r = 4'b0111;
      end
      5'h0a : begin
        color_bar_color_r = 4'b0111;
      end
      5'h0b : begin
        color_bar_color_r = 4'b0111;
      end
      5'h0c : begin
        color_bar_color_r = 4'b1111;
      end
      5'h0d : begin
        color_bar_color_r = 4'b1111;
      end
      5'h0e : begin
        color_bar_color_r = 4'b1111;
      end
      5'h0f : begin
        color_bar_color_r = 4'b1111;
      end
      5'h10 : begin
        color_bar_color_r = 4'b1111;
      end
      5'h11 : begin
        color_bar_color_r = 4'b1111;
      end
      5'h12 : begin
        color_bar_color_r = 4'b1111;
      end
      5'h13 : begin
        color_bar_color_r = 4'b1111;
      end
      default : begin
        color_bar_color_r = 4'b1111;
      end
    endcase
  end

  assign color_palette_idx = {_zz_color_palette_idx,_zz_color_palette_idx_2};
  assign color_palette_color_vec_0 = color_palette_idx[3 : 0];
  assign color_palette_color_vec_1 = color_palette_idx[7 : 4];
  assign color_palette_color_vec_2 = color_palette_idx[11 : 8];
  always @(*) begin
    color_palette_color_r = color_palette_color_vec_2;
    if(when_patgen_l87) begin
      color_palette_color_r[3] = 1'b1;
    end
  end

  assign color_palette_color_g = color_palette_color_vec_1;
  assign color_palette_color_b = color_palette_color_vec_0;
  assign when_patgen_l87 = (sel_id_value == 2'b10);
  always @(*) begin
    case(sel_id_value)
      2'b00 : begin
        _zz_io_color_r = color_bar_color_r;
      end
      2'b01, 2'b10 : begin
        _zz_io_color_r = color_palette_color_r;
      end
      default : begin
        _zz_io_color_r = color_blank_r;
      end
    endcase
  end

  always @(*) begin
    case(sel_id_value)
      2'b00 : begin
        _zz_io_color_g = color_bar_color_g;
      end
      2'b01, 2'b10 : begin
        _zz_io_color_g = color_palette_color_g;
      end
      default : begin
        _zz_io_color_g = color_blank_g;
      end
    endcase
  end

  always @(*) begin
    case(sel_id_value)
      2'b00 : begin
        _zz_io_color_b = color_bar_color_b;
      end
      2'b01, 2'b10 : begin
        _zz_io_color_b = color_palette_color_b;
      end
      default : begin
        _zz_io_color_b = color_blank_b;
      end
    endcase
  end

  assign io_color_r = _zz_io_color_r;
  assign io_color_g = _zz_io_color_g;
  assign io_color_b = _zz_io_color_b;
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      sel_id_value <= 2'b00;
    end else begin
      sel_id_value <= sel_id_valueNext;
    end
  end


endmodule

module layout (
  input      [9:0]    io_x,
  input      [9:0]    io_y,
  output reg          io_inside,
  output     [3:0]    io_color_r,
  output     [3:0]    io_color_g,
  output     [3:0]    io_color_b,
  input               clk,
  input               reset
);

  wire                rectangle_1_io_inside;
  wire       [3:0]    rectangle_1_io_color_r;
  wire       [3:0]    rectangle_1_io_color_g;
  wire       [3:0]    rectangle_1_io_color_b;
  wire                square_1_io_inside;
  wire       [3:0]    square_1_io_color_r;
  wire       [3:0]    square_1_io_color_g;
  wire       [3:0]    square_1_io_color_b;
  wire                ball_1_io_inside;
  wire       [3:0]    ball_1_io_color_r;
  wire       [3:0]    ball_1_io_color_g;
  wire       [3:0]    ball_1_io_color_b;
  reg        [3:0]    color_out_r;
  reg        [3:0]    color_out_g;
  reg        [3:0]    color_out_b;
  wire                inside_out;

  rectangle rectangle_1 (
    .io_x       (io_x[9:0]                  ), //i
    .io_y       (io_y[9:0]                  ), //i
    .io_inside  (rectangle_1_io_inside      ), //o
    .io_color_r (rectangle_1_io_color_r[3:0]), //o
    .io_color_g (rectangle_1_io_color_g[3:0]), //o
    .io_color_b (rectangle_1_io_color_b[3:0]), //o
    .clk        (clk                        ), //i
    .reset      (reset                      )  //i
  );
  square square_1 (
    .io_x       (io_x[9:0]               ), //i
    .io_y       (io_y[9:0]               ), //i
    .io_inside  (square_1_io_inside      ), //o
    .io_color_r (square_1_io_color_r[3:0]), //o
    .io_color_g (square_1_io_color_g[3:0]), //o
    .io_color_b (square_1_io_color_b[3:0]), //o
    .clk        (clk                     ), //i
    .reset      (reset                   )  //i
  );
  ball ball_1 (
    .io_x       (io_x[9:0]             ), //i
    .io_y       (io_y[9:0]             ), //i
    .io_inside  (ball_1_io_inside      ), //o
    .io_color_r (ball_1_io_color_r[3:0]), //o
    .io_color_g (ball_1_io_color_g[3:0]), //o
    .io_color_b (ball_1_io_color_b[3:0]), //o
    .clk        (clk                   ), //i
    .reset      (reset                 )  //i
  );
  always @(*) begin
    color_out_r = 4'b0000;
    if(rectangle_1_io_inside) begin
      color_out_r = rectangle_1_io_color_r;
    end
    if(square_1_io_inside) begin
      color_out_r = square_1_io_color_r;
    end
    if(ball_1_io_inside) begin
      color_out_r = ball_1_io_color_r;
    end
  end

  always @(*) begin
    color_out_g = 4'b0000;
    if(rectangle_1_io_inside) begin
      color_out_g = rectangle_1_io_color_g;
    end
    if(square_1_io_inside) begin
      color_out_g = square_1_io_color_g;
    end
    if(ball_1_io_inside) begin
      color_out_g = ball_1_io_color_g;
    end
  end

  always @(*) begin
    color_out_b = 4'b0000;
    if(rectangle_1_io_inside) begin
      color_out_b = rectangle_1_io_color_b;
    end
    if(square_1_io_inside) begin
      color_out_b = square_1_io_color_b;
    end
    if(ball_1_io_inside) begin
      color_out_b = ball_1_io_color_b;
    end
  end

  assign inside_out = 1'b0;
  assign io_color_r = color_out_r;
  assign io_color_g = color_out_g;
  assign io_color_b = color_out_b;
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      io_inside <= 1'b0;
    end else begin
      io_inside <= (((inside_out || rectangle_1_io_inside) || square_1_io_inside) || ball_1_io_inside);
    end
  end


endmodule

module ball (
  input      [9:0]    io_x,
  input      [9:0]    io_y,
  output reg          io_inside,
  output     [3:0]    io_color_r,
  output     [3:0]    io_color_g,
  output     [3:0]    io_color_b,
  input               clk,
  input               reset
);

  wire       [9:0]    _zz_x_offset;
  wire       [9:0]    _zz_y_offset;
  reg        [99:0]   _zz_xBits;
  wire       [9:0]    _zz_when_shape_l120;
  wire       [9:0]    _zz_when_shape_l120_1;
  wire       [9:0]    x0;
  wire       [9:0]    y0;
  wire       [9:0]    diameter;
  reg        [99:0]   rom_0;
  reg        [99:0]   rom_1;
  reg        [99:0]   rom_2;
  reg        [99:0]   rom_3;
  reg        [99:0]   rom_4;
  reg        [99:0]   rom_5;
  reg        [99:0]   rom_6;
  reg        [99:0]   rom_7;
  reg        [99:0]   rom_8;
  reg        [99:0]   rom_9;
  reg        [99:0]   rom_10;
  reg        [99:0]   rom_11;
  reg        [99:0]   rom_12;
  reg        [99:0]   rom_13;
  reg        [99:0]   rom_14;
  reg        [99:0]   rom_15;
  reg        [99:0]   rom_16;
  reg        [99:0]   rom_17;
  reg        [99:0]   rom_18;
  reg        [99:0]   rom_19;
  reg        [99:0]   rom_20;
  reg        [99:0]   rom_21;
  reg        [99:0]   rom_22;
  reg        [99:0]   rom_23;
  reg        [99:0]   rom_24;
  reg        [99:0]   rom_25;
  reg        [99:0]   rom_26;
  reg        [99:0]   rom_27;
  reg        [99:0]   rom_28;
  reg        [99:0]   rom_29;
  reg        [99:0]   rom_30;
  reg        [99:0]   rom_31;
  reg        [99:0]   rom_32;
  reg        [99:0]   rom_33;
  reg        [99:0]   rom_34;
  reg        [99:0]   rom_35;
  reg        [99:0]   rom_36;
  reg        [99:0]   rom_37;
  reg        [99:0]   rom_38;
  reg        [99:0]   rom_39;
  reg        [99:0]   rom_40;
  reg        [99:0]   rom_41;
  reg        [99:0]   rom_42;
  reg        [99:0]   rom_43;
  reg        [99:0]   rom_44;
  reg        [99:0]   rom_45;
  reg        [99:0]   rom_46;
  reg        [99:0]   rom_47;
  reg        [99:0]   rom_48;
  reg        [99:0]   rom_49;
  reg        [99:0]   rom_50;
  reg        [99:0]   rom_51;
  reg        [99:0]   rom_52;
  reg        [99:0]   rom_53;
  reg        [99:0]   rom_54;
  reg        [99:0]   rom_55;
  reg        [99:0]   rom_56;
  reg        [99:0]   rom_57;
  reg        [99:0]   rom_58;
  reg        [99:0]   rom_59;
  reg        [99:0]   rom_60;
  reg        [99:0]   rom_61;
  reg        [99:0]   rom_62;
  reg        [99:0]   rom_63;
  reg        [99:0]   rom_64;
  reg        [99:0]   rom_65;
  reg        [99:0]   rom_66;
  reg        [99:0]   rom_67;
  reg        [99:0]   rom_68;
  reg        [99:0]   rom_69;
  reg        [99:0]   rom_70;
  reg        [99:0]   rom_71;
  reg        [99:0]   rom_72;
  reg        [99:0]   rom_73;
  reg        [99:0]   rom_74;
  reg        [99:0]   rom_75;
  reg        [99:0]   rom_76;
  reg        [99:0]   rom_77;
  reg        [99:0]   rom_78;
  reg        [99:0]   rom_79;
  reg        [99:0]   rom_80;
  reg        [99:0]   rom_81;
  reg        [99:0]   rom_82;
  reg        [99:0]   rom_83;
  reg        [99:0]   rom_84;
  reg        [99:0]   rom_85;
  reg        [99:0]   rom_86;
  reg        [99:0]   rom_87;
  reg        [99:0]   rom_88;
  reg        [99:0]   rom_89;
  reg        [99:0]   rom_90;
  reg        [99:0]   rom_91;
  reg        [99:0]   rom_92;
  reg        [99:0]   rom_93;
  reg        [99:0]   rom_94;
  reg        [99:0]   rom_95;
  reg        [99:0]   rom_96;
  reg        [99:0]   rom_97;
  reg        [99:0]   rom_98;
  reg        [99:0]   rom_99;
  wire       [6:0]    x_offset;
  wire       [6:0]    y_offset;
  wire       [99:0]   xBits;
  wire                when_shape_l120;
  function [99:0] zz_rom_0(input dummy);
    begin
      zz_rom_0[0] = 1'b0;
      zz_rom_0[1] = 1'b0;
      zz_rom_0[2] = 1'b0;
      zz_rom_0[3] = 1'b0;
      zz_rom_0[4] = 1'b0;
      zz_rom_0[5] = 1'b0;
      zz_rom_0[6] = 1'b0;
      zz_rom_0[7] = 1'b0;
      zz_rom_0[8] = 1'b0;
      zz_rom_0[9] = 1'b0;
      zz_rom_0[10] = 1'b0;
      zz_rom_0[11] = 1'b0;
      zz_rom_0[12] = 1'b0;
      zz_rom_0[13] = 1'b0;
      zz_rom_0[14] = 1'b0;
      zz_rom_0[15] = 1'b0;
      zz_rom_0[16] = 1'b0;
      zz_rom_0[17] = 1'b0;
      zz_rom_0[18] = 1'b0;
      zz_rom_0[19] = 1'b0;
      zz_rom_0[20] = 1'b0;
      zz_rom_0[21] = 1'b0;
      zz_rom_0[22] = 1'b0;
      zz_rom_0[23] = 1'b0;
      zz_rom_0[24] = 1'b0;
      zz_rom_0[25] = 1'b0;
      zz_rom_0[26] = 1'b0;
      zz_rom_0[27] = 1'b0;
      zz_rom_0[28] = 1'b0;
      zz_rom_0[29] = 1'b0;
      zz_rom_0[30] = 1'b0;
      zz_rom_0[31] = 1'b0;
      zz_rom_0[32] = 1'b0;
      zz_rom_0[33] = 1'b0;
      zz_rom_0[34] = 1'b0;
      zz_rom_0[35] = 1'b0;
      zz_rom_0[36] = 1'b0;
      zz_rom_0[37] = 1'b0;
      zz_rom_0[38] = 1'b0;
      zz_rom_0[39] = 1'b0;
      zz_rom_0[40] = 1'b0;
      zz_rom_0[41] = 1'b0;
      zz_rom_0[42] = 1'b0;
      zz_rom_0[43] = 1'b0;
      zz_rom_0[44] = 1'b0;
      zz_rom_0[45] = 1'b0;
      zz_rom_0[46] = 1'b0;
      zz_rom_0[47] = 1'b0;
      zz_rom_0[48] = 1'b0;
      zz_rom_0[49] = 1'b0;
      zz_rom_0[50] = 1'b1;
      zz_rom_0[51] = 1'b0;
      zz_rom_0[52] = 1'b0;
      zz_rom_0[53] = 1'b0;
      zz_rom_0[54] = 1'b0;
      zz_rom_0[55] = 1'b0;
      zz_rom_0[56] = 1'b0;
      zz_rom_0[57] = 1'b0;
      zz_rom_0[58] = 1'b0;
      zz_rom_0[59] = 1'b0;
      zz_rom_0[60] = 1'b0;
      zz_rom_0[61] = 1'b0;
      zz_rom_0[62] = 1'b0;
      zz_rom_0[63] = 1'b0;
      zz_rom_0[64] = 1'b0;
      zz_rom_0[65] = 1'b0;
      zz_rom_0[66] = 1'b0;
      zz_rom_0[67] = 1'b0;
      zz_rom_0[68] = 1'b0;
      zz_rom_0[69] = 1'b0;
      zz_rom_0[70] = 1'b0;
      zz_rom_0[71] = 1'b0;
      zz_rom_0[72] = 1'b0;
      zz_rom_0[73] = 1'b0;
      zz_rom_0[74] = 1'b0;
      zz_rom_0[75] = 1'b0;
      zz_rom_0[76] = 1'b0;
      zz_rom_0[77] = 1'b0;
      zz_rom_0[78] = 1'b0;
      zz_rom_0[79] = 1'b0;
      zz_rom_0[80] = 1'b0;
      zz_rom_0[81] = 1'b0;
      zz_rom_0[82] = 1'b0;
      zz_rom_0[83] = 1'b0;
      zz_rom_0[84] = 1'b0;
      zz_rom_0[85] = 1'b0;
      zz_rom_0[86] = 1'b0;
      zz_rom_0[87] = 1'b0;
      zz_rom_0[88] = 1'b0;
      zz_rom_0[89] = 1'b0;
      zz_rom_0[90] = 1'b0;
      zz_rom_0[91] = 1'b0;
      zz_rom_0[92] = 1'b0;
      zz_rom_0[93] = 1'b0;
      zz_rom_0[94] = 1'b0;
      zz_rom_0[95] = 1'b0;
      zz_rom_0[96] = 1'b0;
      zz_rom_0[97] = 1'b0;
      zz_rom_0[98] = 1'b0;
      zz_rom_0[99] = 1'b0;
    end
  endfunction
  wire [99:0] _zz_1;
  function [99:0] zz_rom_1(input dummy);
    begin
      zz_rom_1[0] = 1'b0;
      zz_rom_1[1] = 1'b0;
      zz_rom_1[2] = 1'b0;
      zz_rom_1[3] = 1'b0;
      zz_rom_1[4] = 1'b0;
      zz_rom_1[5] = 1'b0;
      zz_rom_1[6] = 1'b0;
      zz_rom_1[7] = 1'b0;
      zz_rom_1[8] = 1'b0;
      zz_rom_1[9] = 1'b0;
      zz_rom_1[10] = 1'b0;
      zz_rom_1[11] = 1'b0;
      zz_rom_1[12] = 1'b0;
      zz_rom_1[13] = 1'b0;
      zz_rom_1[14] = 1'b0;
      zz_rom_1[15] = 1'b0;
      zz_rom_1[16] = 1'b0;
      zz_rom_1[17] = 1'b0;
      zz_rom_1[18] = 1'b0;
      zz_rom_1[19] = 1'b0;
      zz_rom_1[20] = 1'b0;
      zz_rom_1[21] = 1'b0;
      zz_rom_1[22] = 1'b0;
      zz_rom_1[23] = 1'b0;
      zz_rom_1[24] = 1'b0;
      zz_rom_1[25] = 1'b0;
      zz_rom_1[26] = 1'b0;
      zz_rom_1[27] = 1'b0;
      zz_rom_1[28] = 1'b0;
      zz_rom_1[29] = 1'b0;
      zz_rom_1[30] = 1'b0;
      zz_rom_1[31] = 1'b0;
      zz_rom_1[32] = 1'b0;
      zz_rom_1[33] = 1'b0;
      zz_rom_1[34] = 1'b0;
      zz_rom_1[35] = 1'b0;
      zz_rom_1[36] = 1'b0;
      zz_rom_1[37] = 1'b0;
      zz_rom_1[38] = 1'b0;
      zz_rom_1[39] = 1'b0;
      zz_rom_1[40] = 1'b0;
      zz_rom_1[41] = 1'b1;
      zz_rom_1[42] = 1'b1;
      zz_rom_1[43] = 1'b1;
      zz_rom_1[44] = 1'b1;
      zz_rom_1[45] = 1'b1;
      zz_rom_1[46] = 1'b1;
      zz_rom_1[47] = 1'b1;
      zz_rom_1[48] = 1'b1;
      zz_rom_1[49] = 1'b1;
      zz_rom_1[50] = 1'b1;
      zz_rom_1[51] = 1'b1;
      zz_rom_1[52] = 1'b1;
      zz_rom_1[53] = 1'b1;
      zz_rom_1[54] = 1'b1;
      zz_rom_1[55] = 1'b1;
      zz_rom_1[56] = 1'b1;
      zz_rom_1[57] = 1'b1;
      zz_rom_1[58] = 1'b1;
      zz_rom_1[59] = 1'b1;
      zz_rom_1[60] = 1'b0;
      zz_rom_1[61] = 1'b0;
      zz_rom_1[62] = 1'b0;
      zz_rom_1[63] = 1'b0;
      zz_rom_1[64] = 1'b0;
      zz_rom_1[65] = 1'b0;
      zz_rom_1[66] = 1'b0;
      zz_rom_1[67] = 1'b0;
      zz_rom_1[68] = 1'b0;
      zz_rom_1[69] = 1'b0;
      zz_rom_1[70] = 1'b0;
      zz_rom_1[71] = 1'b0;
      zz_rom_1[72] = 1'b0;
      zz_rom_1[73] = 1'b0;
      zz_rom_1[74] = 1'b0;
      zz_rom_1[75] = 1'b0;
      zz_rom_1[76] = 1'b0;
      zz_rom_1[77] = 1'b0;
      zz_rom_1[78] = 1'b0;
      zz_rom_1[79] = 1'b0;
      zz_rom_1[80] = 1'b0;
      zz_rom_1[81] = 1'b0;
      zz_rom_1[82] = 1'b0;
      zz_rom_1[83] = 1'b0;
      zz_rom_1[84] = 1'b0;
      zz_rom_1[85] = 1'b0;
      zz_rom_1[86] = 1'b0;
      zz_rom_1[87] = 1'b0;
      zz_rom_1[88] = 1'b0;
      zz_rom_1[89] = 1'b0;
      zz_rom_1[90] = 1'b0;
      zz_rom_1[91] = 1'b0;
      zz_rom_1[92] = 1'b0;
      zz_rom_1[93] = 1'b0;
      zz_rom_1[94] = 1'b0;
      zz_rom_1[95] = 1'b0;
      zz_rom_1[96] = 1'b0;
      zz_rom_1[97] = 1'b0;
      zz_rom_1[98] = 1'b0;
      zz_rom_1[99] = 1'b0;
    end
  endfunction
  wire [99:0] _zz_2;
  function [99:0] zz_rom_2(input dummy);
    begin
      zz_rom_2[0] = 1'b0;
      zz_rom_2[1] = 1'b0;
      zz_rom_2[2] = 1'b0;
      zz_rom_2[3] = 1'b0;
      zz_rom_2[4] = 1'b0;
      zz_rom_2[5] = 1'b0;
      zz_rom_2[6] = 1'b0;
      zz_rom_2[7] = 1'b0;
      zz_rom_2[8] = 1'b0;
      zz_rom_2[9] = 1'b0;
      zz_rom_2[10] = 1'b0;
      zz_rom_2[11] = 1'b0;
      zz_rom_2[12] = 1'b0;
      zz_rom_2[13] = 1'b0;
      zz_rom_2[14] = 1'b0;
      zz_rom_2[15] = 1'b0;
      zz_rom_2[16] = 1'b0;
      zz_rom_2[17] = 1'b0;
      zz_rom_2[18] = 1'b0;
      zz_rom_2[19] = 1'b0;
      zz_rom_2[20] = 1'b0;
      zz_rom_2[21] = 1'b0;
      zz_rom_2[22] = 1'b0;
      zz_rom_2[23] = 1'b0;
      zz_rom_2[24] = 1'b0;
      zz_rom_2[25] = 1'b0;
      zz_rom_2[26] = 1'b0;
      zz_rom_2[27] = 1'b0;
      zz_rom_2[28] = 1'b0;
      zz_rom_2[29] = 1'b0;
      zz_rom_2[30] = 1'b0;
      zz_rom_2[31] = 1'b0;
      zz_rom_2[32] = 1'b0;
      zz_rom_2[33] = 1'b0;
      zz_rom_2[34] = 1'b0;
      zz_rom_2[35] = 1'b0;
      zz_rom_2[36] = 1'b1;
      zz_rom_2[37] = 1'b1;
      zz_rom_2[38] = 1'b1;
      zz_rom_2[39] = 1'b1;
      zz_rom_2[40] = 1'b1;
      zz_rom_2[41] = 1'b1;
      zz_rom_2[42] = 1'b1;
      zz_rom_2[43] = 1'b1;
      zz_rom_2[44] = 1'b1;
      zz_rom_2[45] = 1'b1;
      zz_rom_2[46] = 1'b1;
      zz_rom_2[47] = 1'b1;
      zz_rom_2[48] = 1'b1;
      zz_rom_2[49] = 1'b1;
      zz_rom_2[50] = 1'b1;
      zz_rom_2[51] = 1'b1;
      zz_rom_2[52] = 1'b1;
      zz_rom_2[53] = 1'b1;
      zz_rom_2[54] = 1'b1;
      zz_rom_2[55] = 1'b1;
      zz_rom_2[56] = 1'b1;
      zz_rom_2[57] = 1'b1;
      zz_rom_2[58] = 1'b1;
      zz_rom_2[59] = 1'b1;
      zz_rom_2[60] = 1'b1;
      zz_rom_2[61] = 1'b1;
      zz_rom_2[62] = 1'b1;
      zz_rom_2[63] = 1'b1;
      zz_rom_2[64] = 1'b1;
      zz_rom_2[65] = 1'b0;
      zz_rom_2[66] = 1'b0;
      zz_rom_2[67] = 1'b0;
      zz_rom_2[68] = 1'b0;
      zz_rom_2[69] = 1'b0;
      zz_rom_2[70] = 1'b0;
      zz_rom_2[71] = 1'b0;
      zz_rom_2[72] = 1'b0;
      zz_rom_2[73] = 1'b0;
      zz_rom_2[74] = 1'b0;
      zz_rom_2[75] = 1'b0;
      zz_rom_2[76] = 1'b0;
      zz_rom_2[77] = 1'b0;
      zz_rom_2[78] = 1'b0;
      zz_rom_2[79] = 1'b0;
      zz_rom_2[80] = 1'b0;
      zz_rom_2[81] = 1'b0;
      zz_rom_2[82] = 1'b0;
      zz_rom_2[83] = 1'b0;
      zz_rom_2[84] = 1'b0;
      zz_rom_2[85] = 1'b0;
      zz_rom_2[86] = 1'b0;
      zz_rom_2[87] = 1'b0;
      zz_rom_2[88] = 1'b0;
      zz_rom_2[89] = 1'b0;
      zz_rom_2[90] = 1'b0;
      zz_rom_2[91] = 1'b0;
      zz_rom_2[92] = 1'b0;
      zz_rom_2[93] = 1'b0;
      zz_rom_2[94] = 1'b0;
      zz_rom_2[95] = 1'b0;
      zz_rom_2[96] = 1'b0;
      zz_rom_2[97] = 1'b0;
      zz_rom_2[98] = 1'b0;
      zz_rom_2[99] = 1'b0;
    end
  endfunction
  wire [99:0] _zz_3;
  function [99:0] zz_rom_3(input dummy);
    begin
      zz_rom_3[0] = 1'b0;
      zz_rom_3[1] = 1'b0;
      zz_rom_3[2] = 1'b0;
      zz_rom_3[3] = 1'b0;
      zz_rom_3[4] = 1'b0;
      zz_rom_3[5] = 1'b0;
      zz_rom_3[6] = 1'b0;
      zz_rom_3[7] = 1'b0;
      zz_rom_3[8] = 1'b0;
      zz_rom_3[9] = 1'b0;
      zz_rom_3[10] = 1'b0;
      zz_rom_3[11] = 1'b0;
      zz_rom_3[12] = 1'b0;
      zz_rom_3[13] = 1'b0;
      zz_rom_3[14] = 1'b0;
      zz_rom_3[15] = 1'b0;
      zz_rom_3[16] = 1'b0;
      zz_rom_3[17] = 1'b0;
      zz_rom_3[18] = 1'b0;
      zz_rom_3[19] = 1'b0;
      zz_rom_3[20] = 1'b0;
      zz_rom_3[21] = 1'b0;
      zz_rom_3[22] = 1'b0;
      zz_rom_3[23] = 1'b0;
      zz_rom_3[24] = 1'b0;
      zz_rom_3[25] = 1'b0;
      zz_rom_3[26] = 1'b0;
      zz_rom_3[27] = 1'b0;
      zz_rom_3[28] = 1'b0;
      zz_rom_3[29] = 1'b0;
      zz_rom_3[30] = 1'b0;
      zz_rom_3[31] = 1'b0;
      zz_rom_3[32] = 1'b0;
      zz_rom_3[33] = 1'b1;
      zz_rom_3[34] = 1'b1;
      zz_rom_3[35] = 1'b1;
      zz_rom_3[36] = 1'b1;
      zz_rom_3[37] = 1'b1;
      zz_rom_3[38] = 1'b1;
      zz_rom_3[39] = 1'b1;
      zz_rom_3[40] = 1'b1;
      zz_rom_3[41] = 1'b1;
      zz_rom_3[42] = 1'b1;
      zz_rom_3[43] = 1'b1;
      zz_rom_3[44] = 1'b1;
      zz_rom_3[45] = 1'b1;
      zz_rom_3[46] = 1'b1;
      zz_rom_3[47] = 1'b1;
      zz_rom_3[48] = 1'b1;
      zz_rom_3[49] = 1'b1;
      zz_rom_3[50] = 1'b1;
      zz_rom_3[51] = 1'b1;
      zz_rom_3[52] = 1'b1;
      zz_rom_3[53] = 1'b1;
      zz_rom_3[54] = 1'b1;
      zz_rom_3[55] = 1'b1;
      zz_rom_3[56] = 1'b1;
      zz_rom_3[57] = 1'b1;
      zz_rom_3[58] = 1'b1;
      zz_rom_3[59] = 1'b1;
      zz_rom_3[60] = 1'b1;
      zz_rom_3[61] = 1'b1;
      zz_rom_3[62] = 1'b1;
      zz_rom_3[63] = 1'b1;
      zz_rom_3[64] = 1'b1;
      zz_rom_3[65] = 1'b1;
      zz_rom_3[66] = 1'b1;
      zz_rom_3[67] = 1'b1;
      zz_rom_3[68] = 1'b0;
      zz_rom_3[69] = 1'b0;
      zz_rom_3[70] = 1'b0;
      zz_rom_3[71] = 1'b0;
      zz_rom_3[72] = 1'b0;
      zz_rom_3[73] = 1'b0;
      zz_rom_3[74] = 1'b0;
      zz_rom_3[75] = 1'b0;
      zz_rom_3[76] = 1'b0;
      zz_rom_3[77] = 1'b0;
      zz_rom_3[78] = 1'b0;
      zz_rom_3[79] = 1'b0;
      zz_rom_3[80] = 1'b0;
      zz_rom_3[81] = 1'b0;
      zz_rom_3[82] = 1'b0;
      zz_rom_3[83] = 1'b0;
      zz_rom_3[84] = 1'b0;
      zz_rom_3[85] = 1'b0;
      zz_rom_3[86] = 1'b0;
      zz_rom_3[87] = 1'b0;
      zz_rom_3[88] = 1'b0;
      zz_rom_3[89] = 1'b0;
      zz_rom_3[90] = 1'b0;
      zz_rom_3[91] = 1'b0;
      zz_rom_3[92] = 1'b0;
      zz_rom_3[93] = 1'b0;
      zz_rom_3[94] = 1'b0;
      zz_rom_3[95] = 1'b0;
      zz_rom_3[96] = 1'b0;
      zz_rom_3[97] = 1'b0;
      zz_rom_3[98] = 1'b0;
      zz_rom_3[99] = 1'b0;
    end
  endfunction
  wire [99:0] _zz_4;
  function [99:0] zz_rom_4(input dummy);
    begin
      zz_rom_4[0] = 1'b0;
      zz_rom_4[1] = 1'b0;
      zz_rom_4[2] = 1'b0;
      zz_rom_4[3] = 1'b0;
      zz_rom_4[4] = 1'b0;
      zz_rom_4[5] = 1'b0;
      zz_rom_4[6] = 1'b0;
      zz_rom_4[7] = 1'b0;
      zz_rom_4[8] = 1'b0;
      zz_rom_4[9] = 1'b0;
      zz_rom_4[10] = 1'b0;
      zz_rom_4[11] = 1'b0;
      zz_rom_4[12] = 1'b0;
      zz_rom_4[13] = 1'b0;
      zz_rom_4[14] = 1'b0;
      zz_rom_4[15] = 1'b0;
      zz_rom_4[16] = 1'b0;
      zz_rom_4[17] = 1'b0;
      zz_rom_4[18] = 1'b0;
      zz_rom_4[19] = 1'b0;
      zz_rom_4[20] = 1'b0;
      zz_rom_4[21] = 1'b0;
      zz_rom_4[22] = 1'b0;
      zz_rom_4[23] = 1'b0;
      zz_rom_4[24] = 1'b0;
      zz_rom_4[25] = 1'b0;
      zz_rom_4[26] = 1'b0;
      zz_rom_4[27] = 1'b0;
      zz_rom_4[28] = 1'b0;
      zz_rom_4[29] = 1'b0;
      zz_rom_4[30] = 1'b0;
      zz_rom_4[31] = 1'b1;
      zz_rom_4[32] = 1'b1;
      zz_rom_4[33] = 1'b1;
      zz_rom_4[34] = 1'b1;
      zz_rom_4[35] = 1'b1;
      zz_rom_4[36] = 1'b1;
      zz_rom_4[37] = 1'b1;
      zz_rom_4[38] = 1'b1;
      zz_rom_4[39] = 1'b1;
      zz_rom_4[40] = 1'b1;
      zz_rom_4[41] = 1'b1;
      zz_rom_4[42] = 1'b1;
      zz_rom_4[43] = 1'b1;
      zz_rom_4[44] = 1'b1;
      zz_rom_4[45] = 1'b1;
      zz_rom_4[46] = 1'b1;
      zz_rom_4[47] = 1'b1;
      zz_rom_4[48] = 1'b1;
      zz_rom_4[49] = 1'b1;
      zz_rom_4[50] = 1'b1;
      zz_rom_4[51] = 1'b1;
      zz_rom_4[52] = 1'b1;
      zz_rom_4[53] = 1'b1;
      zz_rom_4[54] = 1'b1;
      zz_rom_4[55] = 1'b1;
      zz_rom_4[56] = 1'b1;
      zz_rom_4[57] = 1'b1;
      zz_rom_4[58] = 1'b1;
      zz_rom_4[59] = 1'b1;
      zz_rom_4[60] = 1'b1;
      zz_rom_4[61] = 1'b1;
      zz_rom_4[62] = 1'b1;
      zz_rom_4[63] = 1'b1;
      zz_rom_4[64] = 1'b1;
      zz_rom_4[65] = 1'b1;
      zz_rom_4[66] = 1'b1;
      zz_rom_4[67] = 1'b1;
      zz_rom_4[68] = 1'b1;
      zz_rom_4[69] = 1'b1;
      zz_rom_4[70] = 1'b0;
      zz_rom_4[71] = 1'b0;
      zz_rom_4[72] = 1'b0;
      zz_rom_4[73] = 1'b0;
      zz_rom_4[74] = 1'b0;
      zz_rom_4[75] = 1'b0;
      zz_rom_4[76] = 1'b0;
      zz_rom_4[77] = 1'b0;
      zz_rom_4[78] = 1'b0;
      zz_rom_4[79] = 1'b0;
      zz_rom_4[80] = 1'b0;
      zz_rom_4[81] = 1'b0;
      zz_rom_4[82] = 1'b0;
      zz_rom_4[83] = 1'b0;
      zz_rom_4[84] = 1'b0;
      zz_rom_4[85] = 1'b0;
      zz_rom_4[86] = 1'b0;
      zz_rom_4[87] = 1'b0;
      zz_rom_4[88] = 1'b0;
      zz_rom_4[89] = 1'b0;
      zz_rom_4[90] = 1'b0;
      zz_rom_4[91] = 1'b0;
      zz_rom_4[92] = 1'b0;
      zz_rom_4[93] = 1'b0;
      zz_rom_4[94] = 1'b0;
      zz_rom_4[95] = 1'b0;
      zz_rom_4[96] = 1'b0;
      zz_rom_4[97] = 1'b0;
      zz_rom_4[98] = 1'b0;
      zz_rom_4[99] = 1'b0;
    end
  endfunction
  wire [99:0] _zz_5;
  function [99:0] zz_rom_5(input dummy);
    begin
      zz_rom_5[0] = 1'b0;
      zz_rom_5[1] = 1'b0;
      zz_rom_5[2] = 1'b0;
      zz_rom_5[3] = 1'b0;
      zz_rom_5[4] = 1'b0;
      zz_rom_5[5] = 1'b0;
      zz_rom_5[6] = 1'b0;
      zz_rom_5[7] = 1'b0;
      zz_rom_5[8] = 1'b0;
      zz_rom_5[9] = 1'b0;
      zz_rom_5[10] = 1'b0;
      zz_rom_5[11] = 1'b0;
      zz_rom_5[12] = 1'b0;
      zz_rom_5[13] = 1'b0;
      zz_rom_5[14] = 1'b0;
      zz_rom_5[15] = 1'b0;
      zz_rom_5[16] = 1'b0;
      zz_rom_5[17] = 1'b0;
      zz_rom_5[18] = 1'b0;
      zz_rom_5[19] = 1'b0;
      zz_rom_5[20] = 1'b0;
      zz_rom_5[21] = 1'b0;
      zz_rom_5[22] = 1'b0;
      zz_rom_5[23] = 1'b0;
      zz_rom_5[24] = 1'b0;
      zz_rom_5[25] = 1'b0;
      zz_rom_5[26] = 1'b0;
      zz_rom_5[27] = 1'b0;
      zz_rom_5[28] = 1'b0;
      zz_rom_5[29] = 1'b1;
      zz_rom_5[30] = 1'b1;
      zz_rom_5[31] = 1'b1;
      zz_rom_5[32] = 1'b1;
      zz_rom_5[33] = 1'b1;
      zz_rom_5[34] = 1'b1;
      zz_rom_5[35] = 1'b1;
      zz_rom_5[36] = 1'b1;
      zz_rom_5[37] = 1'b1;
      zz_rom_5[38] = 1'b1;
      zz_rom_5[39] = 1'b1;
      zz_rom_5[40] = 1'b1;
      zz_rom_5[41] = 1'b1;
      zz_rom_5[42] = 1'b1;
      zz_rom_5[43] = 1'b1;
      zz_rom_5[44] = 1'b1;
      zz_rom_5[45] = 1'b1;
      zz_rom_5[46] = 1'b1;
      zz_rom_5[47] = 1'b1;
      zz_rom_5[48] = 1'b1;
      zz_rom_5[49] = 1'b1;
      zz_rom_5[50] = 1'b1;
      zz_rom_5[51] = 1'b1;
      zz_rom_5[52] = 1'b1;
      zz_rom_5[53] = 1'b1;
      zz_rom_5[54] = 1'b1;
      zz_rom_5[55] = 1'b1;
      zz_rom_5[56] = 1'b1;
      zz_rom_5[57] = 1'b1;
      zz_rom_5[58] = 1'b1;
      zz_rom_5[59] = 1'b1;
      zz_rom_5[60] = 1'b1;
      zz_rom_5[61] = 1'b1;
      zz_rom_5[62] = 1'b1;
      zz_rom_5[63] = 1'b1;
      zz_rom_5[64] = 1'b1;
      zz_rom_5[65] = 1'b1;
      zz_rom_5[66] = 1'b1;
      zz_rom_5[67] = 1'b1;
      zz_rom_5[68] = 1'b1;
      zz_rom_5[69] = 1'b1;
      zz_rom_5[70] = 1'b1;
      zz_rom_5[71] = 1'b1;
      zz_rom_5[72] = 1'b0;
      zz_rom_5[73] = 1'b0;
      zz_rom_5[74] = 1'b0;
      zz_rom_5[75] = 1'b0;
      zz_rom_5[76] = 1'b0;
      zz_rom_5[77] = 1'b0;
      zz_rom_5[78] = 1'b0;
      zz_rom_5[79] = 1'b0;
      zz_rom_5[80] = 1'b0;
      zz_rom_5[81] = 1'b0;
      zz_rom_5[82] = 1'b0;
      zz_rom_5[83] = 1'b0;
      zz_rom_5[84] = 1'b0;
      zz_rom_5[85] = 1'b0;
      zz_rom_5[86] = 1'b0;
      zz_rom_5[87] = 1'b0;
      zz_rom_5[88] = 1'b0;
      zz_rom_5[89] = 1'b0;
      zz_rom_5[90] = 1'b0;
      zz_rom_5[91] = 1'b0;
      zz_rom_5[92] = 1'b0;
      zz_rom_5[93] = 1'b0;
      zz_rom_5[94] = 1'b0;
      zz_rom_5[95] = 1'b0;
      zz_rom_5[96] = 1'b0;
      zz_rom_5[97] = 1'b0;
      zz_rom_5[98] = 1'b0;
      zz_rom_5[99] = 1'b0;
    end
  endfunction
  wire [99:0] _zz_6;
  function [99:0] zz_rom_6(input dummy);
    begin
      zz_rom_6[0] = 1'b0;
      zz_rom_6[1] = 1'b0;
      zz_rom_6[2] = 1'b0;
      zz_rom_6[3] = 1'b0;
      zz_rom_6[4] = 1'b0;
      zz_rom_6[5] = 1'b0;
      zz_rom_6[6] = 1'b0;
      zz_rom_6[7] = 1'b0;
      zz_rom_6[8] = 1'b0;
      zz_rom_6[9] = 1'b0;
      zz_rom_6[10] = 1'b0;
      zz_rom_6[11] = 1'b0;
      zz_rom_6[12] = 1'b0;
      zz_rom_6[13] = 1'b0;
      zz_rom_6[14] = 1'b0;
      zz_rom_6[15] = 1'b0;
      zz_rom_6[16] = 1'b0;
      zz_rom_6[17] = 1'b0;
      zz_rom_6[18] = 1'b0;
      zz_rom_6[19] = 1'b0;
      zz_rom_6[20] = 1'b0;
      zz_rom_6[21] = 1'b0;
      zz_rom_6[22] = 1'b0;
      zz_rom_6[23] = 1'b0;
      zz_rom_6[24] = 1'b0;
      zz_rom_6[25] = 1'b0;
      zz_rom_6[26] = 1'b0;
      zz_rom_6[27] = 1'b1;
      zz_rom_6[28] = 1'b1;
      zz_rom_6[29] = 1'b1;
      zz_rom_6[30] = 1'b1;
      zz_rom_6[31] = 1'b1;
      zz_rom_6[32] = 1'b1;
      zz_rom_6[33] = 1'b1;
      zz_rom_6[34] = 1'b1;
      zz_rom_6[35] = 1'b1;
      zz_rom_6[36] = 1'b1;
      zz_rom_6[37] = 1'b1;
      zz_rom_6[38] = 1'b1;
      zz_rom_6[39] = 1'b1;
      zz_rom_6[40] = 1'b1;
      zz_rom_6[41] = 1'b1;
      zz_rom_6[42] = 1'b1;
      zz_rom_6[43] = 1'b1;
      zz_rom_6[44] = 1'b1;
      zz_rom_6[45] = 1'b1;
      zz_rom_6[46] = 1'b1;
      zz_rom_6[47] = 1'b1;
      zz_rom_6[48] = 1'b1;
      zz_rom_6[49] = 1'b1;
      zz_rom_6[50] = 1'b1;
      zz_rom_6[51] = 1'b1;
      zz_rom_6[52] = 1'b1;
      zz_rom_6[53] = 1'b1;
      zz_rom_6[54] = 1'b1;
      zz_rom_6[55] = 1'b1;
      zz_rom_6[56] = 1'b1;
      zz_rom_6[57] = 1'b1;
      zz_rom_6[58] = 1'b1;
      zz_rom_6[59] = 1'b1;
      zz_rom_6[60] = 1'b1;
      zz_rom_6[61] = 1'b1;
      zz_rom_6[62] = 1'b1;
      zz_rom_6[63] = 1'b1;
      zz_rom_6[64] = 1'b1;
      zz_rom_6[65] = 1'b1;
      zz_rom_6[66] = 1'b1;
      zz_rom_6[67] = 1'b1;
      zz_rom_6[68] = 1'b1;
      zz_rom_6[69] = 1'b1;
      zz_rom_6[70] = 1'b1;
      zz_rom_6[71] = 1'b1;
      zz_rom_6[72] = 1'b1;
      zz_rom_6[73] = 1'b1;
      zz_rom_6[74] = 1'b0;
      zz_rom_6[75] = 1'b0;
      zz_rom_6[76] = 1'b0;
      zz_rom_6[77] = 1'b0;
      zz_rom_6[78] = 1'b0;
      zz_rom_6[79] = 1'b0;
      zz_rom_6[80] = 1'b0;
      zz_rom_6[81] = 1'b0;
      zz_rom_6[82] = 1'b0;
      zz_rom_6[83] = 1'b0;
      zz_rom_6[84] = 1'b0;
      zz_rom_6[85] = 1'b0;
      zz_rom_6[86] = 1'b0;
      zz_rom_6[87] = 1'b0;
      zz_rom_6[88] = 1'b0;
      zz_rom_6[89] = 1'b0;
      zz_rom_6[90] = 1'b0;
      zz_rom_6[91] = 1'b0;
      zz_rom_6[92] = 1'b0;
      zz_rom_6[93] = 1'b0;
      zz_rom_6[94] = 1'b0;
      zz_rom_6[95] = 1'b0;
      zz_rom_6[96] = 1'b0;
      zz_rom_6[97] = 1'b0;
      zz_rom_6[98] = 1'b0;
      zz_rom_6[99] = 1'b0;
    end
  endfunction
  wire [99:0] _zz_7;
  function [99:0] zz_rom_7(input dummy);
    begin
      zz_rom_7[0] = 1'b0;
      zz_rom_7[1] = 1'b0;
      zz_rom_7[2] = 1'b0;
      zz_rom_7[3] = 1'b0;
      zz_rom_7[4] = 1'b0;
      zz_rom_7[5] = 1'b0;
      zz_rom_7[6] = 1'b0;
      zz_rom_7[7] = 1'b0;
      zz_rom_7[8] = 1'b0;
      zz_rom_7[9] = 1'b0;
      zz_rom_7[10] = 1'b0;
      zz_rom_7[11] = 1'b0;
      zz_rom_7[12] = 1'b0;
      zz_rom_7[13] = 1'b0;
      zz_rom_7[14] = 1'b0;
      zz_rom_7[15] = 1'b0;
      zz_rom_7[16] = 1'b0;
      zz_rom_7[17] = 1'b0;
      zz_rom_7[18] = 1'b0;
      zz_rom_7[19] = 1'b0;
      zz_rom_7[20] = 1'b0;
      zz_rom_7[21] = 1'b0;
      zz_rom_7[22] = 1'b0;
      zz_rom_7[23] = 1'b0;
      zz_rom_7[24] = 1'b0;
      zz_rom_7[25] = 1'b1;
      zz_rom_7[26] = 1'b1;
      zz_rom_7[27] = 1'b1;
      zz_rom_7[28] = 1'b1;
      zz_rom_7[29] = 1'b1;
      zz_rom_7[30] = 1'b1;
      zz_rom_7[31] = 1'b1;
      zz_rom_7[32] = 1'b1;
      zz_rom_7[33] = 1'b1;
      zz_rom_7[34] = 1'b1;
      zz_rom_7[35] = 1'b1;
      zz_rom_7[36] = 1'b1;
      zz_rom_7[37] = 1'b1;
      zz_rom_7[38] = 1'b1;
      zz_rom_7[39] = 1'b1;
      zz_rom_7[40] = 1'b1;
      zz_rom_7[41] = 1'b1;
      zz_rom_7[42] = 1'b1;
      zz_rom_7[43] = 1'b1;
      zz_rom_7[44] = 1'b1;
      zz_rom_7[45] = 1'b1;
      zz_rom_7[46] = 1'b1;
      zz_rom_7[47] = 1'b1;
      zz_rom_7[48] = 1'b1;
      zz_rom_7[49] = 1'b1;
      zz_rom_7[50] = 1'b1;
      zz_rom_7[51] = 1'b1;
      zz_rom_7[52] = 1'b1;
      zz_rom_7[53] = 1'b1;
      zz_rom_7[54] = 1'b1;
      zz_rom_7[55] = 1'b1;
      zz_rom_7[56] = 1'b1;
      zz_rom_7[57] = 1'b1;
      zz_rom_7[58] = 1'b1;
      zz_rom_7[59] = 1'b1;
      zz_rom_7[60] = 1'b1;
      zz_rom_7[61] = 1'b1;
      zz_rom_7[62] = 1'b1;
      zz_rom_7[63] = 1'b1;
      zz_rom_7[64] = 1'b1;
      zz_rom_7[65] = 1'b1;
      zz_rom_7[66] = 1'b1;
      zz_rom_7[67] = 1'b1;
      zz_rom_7[68] = 1'b1;
      zz_rom_7[69] = 1'b1;
      zz_rom_7[70] = 1'b1;
      zz_rom_7[71] = 1'b1;
      zz_rom_7[72] = 1'b1;
      zz_rom_7[73] = 1'b1;
      zz_rom_7[74] = 1'b1;
      zz_rom_7[75] = 1'b1;
      zz_rom_7[76] = 1'b0;
      zz_rom_7[77] = 1'b0;
      zz_rom_7[78] = 1'b0;
      zz_rom_7[79] = 1'b0;
      zz_rom_7[80] = 1'b0;
      zz_rom_7[81] = 1'b0;
      zz_rom_7[82] = 1'b0;
      zz_rom_7[83] = 1'b0;
      zz_rom_7[84] = 1'b0;
      zz_rom_7[85] = 1'b0;
      zz_rom_7[86] = 1'b0;
      zz_rom_7[87] = 1'b0;
      zz_rom_7[88] = 1'b0;
      zz_rom_7[89] = 1'b0;
      zz_rom_7[90] = 1'b0;
      zz_rom_7[91] = 1'b0;
      zz_rom_7[92] = 1'b0;
      zz_rom_7[93] = 1'b0;
      zz_rom_7[94] = 1'b0;
      zz_rom_7[95] = 1'b0;
      zz_rom_7[96] = 1'b0;
      zz_rom_7[97] = 1'b0;
      zz_rom_7[98] = 1'b0;
      zz_rom_7[99] = 1'b0;
    end
  endfunction
  wire [99:0] _zz_8;
  function [99:0] zz_rom_8(input dummy);
    begin
      zz_rom_8[0] = 1'b0;
      zz_rom_8[1] = 1'b0;
      zz_rom_8[2] = 1'b0;
      zz_rom_8[3] = 1'b0;
      zz_rom_8[4] = 1'b0;
      zz_rom_8[5] = 1'b0;
      zz_rom_8[6] = 1'b0;
      zz_rom_8[7] = 1'b0;
      zz_rom_8[8] = 1'b0;
      zz_rom_8[9] = 1'b0;
      zz_rom_8[10] = 1'b0;
      zz_rom_8[11] = 1'b0;
      zz_rom_8[12] = 1'b0;
      zz_rom_8[13] = 1'b0;
      zz_rom_8[14] = 1'b0;
      zz_rom_8[15] = 1'b0;
      zz_rom_8[16] = 1'b0;
      zz_rom_8[17] = 1'b0;
      zz_rom_8[18] = 1'b0;
      zz_rom_8[19] = 1'b0;
      zz_rom_8[20] = 1'b0;
      zz_rom_8[21] = 1'b0;
      zz_rom_8[22] = 1'b0;
      zz_rom_8[23] = 1'b1;
      zz_rom_8[24] = 1'b1;
      zz_rom_8[25] = 1'b1;
      zz_rom_8[26] = 1'b1;
      zz_rom_8[27] = 1'b1;
      zz_rom_8[28] = 1'b1;
      zz_rom_8[29] = 1'b1;
      zz_rom_8[30] = 1'b1;
      zz_rom_8[31] = 1'b1;
      zz_rom_8[32] = 1'b1;
      zz_rom_8[33] = 1'b1;
      zz_rom_8[34] = 1'b1;
      zz_rom_8[35] = 1'b1;
      zz_rom_8[36] = 1'b1;
      zz_rom_8[37] = 1'b1;
      zz_rom_8[38] = 1'b1;
      zz_rom_8[39] = 1'b1;
      zz_rom_8[40] = 1'b1;
      zz_rom_8[41] = 1'b1;
      zz_rom_8[42] = 1'b1;
      zz_rom_8[43] = 1'b1;
      zz_rom_8[44] = 1'b1;
      zz_rom_8[45] = 1'b1;
      zz_rom_8[46] = 1'b1;
      zz_rom_8[47] = 1'b1;
      zz_rom_8[48] = 1'b1;
      zz_rom_8[49] = 1'b1;
      zz_rom_8[50] = 1'b1;
      zz_rom_8[51] = 1'b1;
      zz_rom_8[52] = 1'b1;
      zz_rom_8[53] = 1'b1;
      zz_rom_8[54] = 1'b1;
      zz_rom_8[55] = 1'b1;
      zz_rom_8[56] = 1'b1;
      zz_rom_8[57] = 1'b1;
      zz_rom_8[58] = 1'b1;
      zz_rom_8[59] = 1'b1;
      zz_rom_8[60] = 1'b1;
      zz_rom_8[61] = 1'b1;
      zz_rom_8[62] = 1'b1;
      zz_rom_8[63] = 1'b1;
      zz_rom_8[64] = 1'b1;
      zz_rom_8[65] = 1'b1;
      zz_rom_8[66] = 1'b1;
      zz_rom_8[67] = 1'b1;
      zz_rom_8[68] = 1'b1;
      zz_rom_8[69] = 1'b1;
      zz_rom_8[70] = 1'b1;
      zz_rom_8[71] = 1'b1;
      zz_rom_8[72] = 1'b1;
      zz_rom_8[73] = 1'b1;
      zz_rom_8[74] = 1'b1;
      zz_rom_8[75] = 1'b1;
      zz_rom_8[76] = 1'b1;
      zz_rom_8[77] = 1'b1;
      zz_rom_8[78] = 1'b0;
      zz_rom_8[79] = 1'b0;
      zz_rom_8[80] = 1'b0;
      zz_rom_8[81] = 1'b0;
      zz_rom_8[82] = 1'b0;
      zz_rom_8[83] = 1'b0;
      zz_rom_8[84] = 1'b0;
      zz_rom_8[85] = 1'b0;
      zz_rom_8[86] = 1'b0;
      zz_rom_8[87] = 1'b0;
      zz_rom_8[88] = 1'b0;
      zz_rom_8[89] = 1'b0;
      zz_rom_8[90] = 1'b0;
      zz_rom_8[91] = 1'b0;
      zz_rom_8[92] = 1'b0;
      zz_rom_8[93] = 1'b0;
      zz_rom_8[94] = 1'b0;
      zz_rom_8[95] = 1'b0;
      zz_rom_8[96] = 1'b0;
      zz_rom_8[97] = 1'b0;
      zz_rom_8[98] = 1'b0;
      zz_rom_8[99] = 1'b0;
    end
  endfunction
  wire [99:0] _zz_9;
  function [99:0] zz_rom_9(input dummy);
    begin
      zz_rom_9[0] = 1'b0;
      zz_rom_9[1] = 1'b0;
      zz_rom_9[2] = 1'b0;
      zz_rom_9[3] = 1'b0;
      zz_rom_9[4] = 1'b0;
      zz_rom_9[5] = 1'b0;
      zz_rom_9[6] = 1'b0;
      zz_rom_9[7] = 1'b0;
      zz_rom_9[8] = 1'b0;
      zz_rom_9[9] = 1'b0;
      zz_rom_9[10] = 1'b0;
      zz_rom_9[11] = 1'b0;
      zz_rom_9[12] = 1'b0;
      zz_rom_9[13] = 1'b0;
      zz_rom_9[14] = 1'b0;
      zz_rom_9[15] = 1'b0;
      zz_rom_9[16] = 1'b0;
      zz_rom_9[17] = 1'b0;
      zz_rom_9[18] = 1'b0;
      zz_rom_9[19] = 1'b0;
      zz_rom_9[20] = 1'b0;
      zz_rom_9[21] = 1'b0;
      zz_rom_9[22] = 1'b1;
      zz_rom_9[23] = 1'b1;
      zz_rom_9[24] = 1'b1;
      zz_rom_9[25] = 1'b1;
      zz_rom_9[26] = 1'b1;
      zz_rom_9[27] = 1'b1;
      zz_rom_9[28] = 1'b1;
      zz_rom_9[29] = 1'b1;
      zz_rom_9[30] = 1'b1;
      zz_rom_9[31] = 1'b1;
      zz_rom_9[32] = 1'b1;
      zz_rom_9[33] = 1'b1;
      zz_rom_9[34] = 1'b1;
      zz_rom_9[35] = 1'b1;
      zz_rom_9[36] = 1'b1;
      zz_rom_9[37] = 1'b1;
      zz_rom_9[38] = 1'b1;
      zz_rom_9[39] = 1'b1;
      zz_rom_9[40] = 1'b1;
      zz_rom_9[41] = 1'b1;
      zz_rom_9[42] = 1'b1;
      zz_rom_9[43] = 1'b1;
      zz_rom_9[44] = 1'b1;
      zz_rom_9[45] = 1'b1;
      zz_rom_9[46] = 1'b1;
      zz_rom_9[47] = 1'b1;
      zz_rom_9[48] = 1'b1;
      zz_rom_9[49] = 1'b1;
      zz_rom_9[50] = 1'b1;
      zz_rom_9[51] = 1'b1;
      zz_rom_9[52] = 1'b1;
      zz_rom_9[53] = 1'b1;
      zz_rom_9[54] = 1'b1;
      zz_rom_9[55] = 1'b1;
      zz_rom_9[56] = 1'b1;
      zz_rom_9[57] = 1'b1;
      zz_rom_9[58] = 1'b1;
      zz_rom_9[59] = 1'b1;
      zz_rom_9[60] = 1'b1;
      zz_rom_9[61] = 1'b1;
      zz_rom_9[62] = 1'b1;
      zz_rom_9[63] = 1'b1;
      zz_rom_9[64] = 1'b1;
      zz_rom_9[65] = 1'b1;
      zz_rom_9[66] = 1'b1;
      zz_rom_9[67] = 1'b1;
      zz_rom_9[68] = 1'b1;
      zz_rom_9[69] = 1'b1;
      zz_rom_9[70] = 1'b1;
      zz_rom_9[71] = 1'b1;
      zz_rom_9[72] = 1'b1;
      zz_rom_9[73] = 1'b1;
      zz_rom_9[74] = 1'b1;
      zz_rom_9[75] = 1'b1;
      zz_rom_9[76] = 1'b1;
      zz_rom_9[77] = 1'b1;
      zz_rom_9[78] = 1'b1;
      zz_rom_9[79] = 1'b0;
      zz_rom_9[80] = 1'b0;
      zz_rom_9[81] = 1'b0;
      zz_rom_9[82] = 1'b0;
      zz_rom_9[83] = 1'b0;
      zz_rom_9[84] = 1'b0;
      zz_rom_9[85] = 1'b0;
      zz_rom_9[86] = 1'b0;
      zz_rom_9[87] = 1'b0;
      zz_rom_9[88] = 1'b0;
      zz_rom_9[89] = 1'b0;
      zz_rom_9[90] = 1'b0;
      zz_rom_9[91] = 1'b0;
      zz_rom_9[92] = 1'b0;
      zz_rom_9[93] = 1'b0;
      zz_rom_9[94] = 1'b0;
      zz_rom_9[95] = 1'b0;
      zz_rom_9[96] = 1'b0;
      zz_rom_9[97] = 1'b0;
      zz_rom_9[98] = 1'b0;
      zz_rom_9[99] = 1'b0;
    end
  endfunction
  wire [99:0] _zz_10;
  function [99:0] zz_rom_10(input dummy);
    begin
      zz_rom_10[0] = 1'b0;
      zz_rom_10[1] = 1'b0;
      zz_rom_10[2] = 1'b0;
      zz_rom_10[3] = 1'b0;
      zz_rom_10[4] = 1'b0;
      zz_rom_10[5] = 1'b0;
      zz_rom_10[6] = 1'b0;
      zz_rom_10[7] = 1'b0;
      zz_rom_10[8] = 1'b0;
      zz_rom_10[9] = 1'b0;
      zz_rom_10[10] = 1'b0;
      zz_rom_10[11] = 1'b0;
      zz_rom_10[12] = 1'b0;
      zz_rom_10[13] = 1'b0;
      zz_rom_10[14] = 1'b0;
      zz_rom_10[15] = 1'b0;
      zz_rom_10[16] = 1'b0;
      zz_rom_10[17] = 1'b0;
      zz_rom_10[18] = 1'b0;
      zz_rom_10[19] = 1'b0;
      zz_rom_10[20] = 1'b1;
      zz_rom_10[21] = 1'b1;
      zz_rom_10[22] = 1'b1;
      zz_rom_10[23] = 1'b1;
      zz_rom_10[24] = 1'b1;
      zz_rom_10[25] = 1'b1;
      zz_rom_10[26] = 1'b1;
      zz_rom_10[27] = 1'b1;
      zz_rom_10[28] = 1'b1;
      zz_rom_10[29] = 1'b1;
      zz_rom_10[30] = 1'b1;
      zz_rom_10[31] = 1'b1;
      zz_rom_10[32] = 1'b1;
      zz_rom_10[33] = 1'b1;
      zz_rom_10[34] = 1'b1;
      zz_rom_10[35] = 1'b1;
      zz_rom_10[36] = 1'b1;
      zz_rom_10[37] = 1'b1;
      zz_rom_10[38] = 1'b1;
      zz_rom_10[39] = 1'b1;
      zz_rom_10[40] = 1'b1;
      zz_rom_10[41] = 1'b1;
      zz_rom_10[42] = 1'b1;
      zz_rom_10[43] = 1'b1;
      zz_rom_10[44] = 1'b1;
      zz_rom_10[45] = 1'b1;
      zz_rom_10[46] = 1'b1;
      zz_rom_10[47] = 1'b1;
      zz_rom_10[48] = 1'b1;
      zz_rom_10[49] = 1'b1;
      zz_rom_10[50] = 1'b1;
      zz_rom_10[51] = 1'b1;
      zz_rom_10[52] = 1'b1;
      zz_rom_10[53] = 1'b1;
      zz_rom_10[54] = 1'b1;
      zz_rom_10[55] = 1'b1;
      zz_rom_10[56] = 1'b1;
      zz_rom_10[57] = 1'b1;
      zz_rom_10[58] = 1'b1;
      zz_rom_10[59] = 1'b1;
      zz_rom_10[60] = 1'b1;
      zz_rom_10[61] = 1'b1;
      zz_rom_10[62] = 1'b1;
      zz_rom_10[63] = 1'b1;
      zz_rom_10[64] = 1'b1;
      zz_rom_10[65] = 1'b1;
      zz_rom_10[66] = 1'b1;
      zz_rom_10[67] = 1'b1;
      zz_rom_10[68] = 1'b1;
      zz_rom_10[69] = 1'b1;
      zz_rom_10[70] = 1'b1;
      zz_rom_10[71] = 1'b1;
      zz_rom_10[72] = 1'b1;
      zz_rom_10[73] = 1'b1;
      zz_rom_10[74] = 1'b1;
      zz_rom_10[75] = 1'b1;
      zz_rom_10[76] = 1'b1;
      zz_rom_10[77] = 1'b1;
      zz_rom_10[78] = 1'b1;
      zz_rom_10[79] = 1'b1;
      zz_rom_10[80] = 1'b1;
      zz_rom_10[81] = 1'b0;
      zz_rom_10[82] = 1'b0;
      zz_rom_10[83] = 1'b0;
      zz_rom_10[84] = 1'b0;
      zz_rom_10[85] = 1'b0;
      zz_rom_10[86] = 1'b0;
      zz_rom_10[87] = 1'b0;
      zz_rom_10[88] = 1'b0;
      zz_rom_10[89] = 1'b0;
      zz_rom_10[90] = 1'b0;
      zz_rom_10[91] = 1'b0;
      zz_rom_10[92] = 1'b0;
      zz_rom_10[93] = 1'b0;
      zz_rom_10[94] = 1'b0;
      zz_rom_10[95] = 1'b0;
      zz_rom_10[96] = 1'b0;
      zz_rom_10[97] = 1'b0;
      zz_rom_10[98] = 1'b0;
      zz_rom_10[99] = 1'b0;
    end
  endfunction
  wire [99:0] _zz_11;
  function [99:0] zz_rom_11(input dummy);
    begin
      zz_rom_11[0] = 1'b0;
      zz_rom_11[1] = 1'b0;
      zz_rom_11[2] = 1'b0;
      zz_rom_11[3] = 1'b0;
      zz_rom_11[4] = 1'b0;
      zz_rom_11[5] = 1'b0;
      zz_rom_11[6] = 1'b0;
      zz_rom_11[7] = 1'b0;
      zz_rom_11[8] = 1'b0;
      zz_rom_11[9] = 1'b0;
      zz_rom_11[10] = 1'b0;
      zz_rom_11[11] = 1'b0;
      zz_rom_11[12] = 1'b0;
      zz_rom_11[13] = 1'b0;
      zz_rom_11[14] = 1'b0;
      zz_rom_11[15] = 1'b0;
      zz_rom_11[16] = 1'b0;
      zz_rom_11[17] = 1'b0;
      zz_rom_11[18] = 1'b0;
      zz_rom_11[19] = 1'b1;
      zz_rom_11[20] = 1'b1;
      zz_rom_11[21] = 1'b1;
      zz_rom_11[22] = 1'b1;
      zz_rom_11[23] = 1'b1;
      zz_rom_11[24] = 1'b1;
      zz_rom_11[25] = 1'b1;
      zz_rom_11[26] = 1'b1;
      zz_rom_11[27] = 1'b1;
      zz_rom_11[28] = 1'b1;
      zz_rom_11[29] = 1'b1;
      zz_rom_11[30] = 1'b1;
      zz_rom_11[31] = 1'b1;
      zz_rom_11[32] = 1'b1;
      zz_rom_11[33] = 1'b1;
      zz_rom_11[34] = 1'b1;
      zz_rom_11[35] = 1'b1;
      zz_rom_11[36] = 1'b1;
      zz_rom_11[37] = 1'b1;
      zz_rom_11[38] = 1'b1;
      zz_rom_11[39] = 1'b1;
      zz_rom_11[40] = 1'b1;
      zz_rom_11[41] = 1'b1;
      zz_rom_11[42] = 1'b1;
      zz_rom_11[43] = 1'b1;
      zz_rom_11[44] = 1'b1;
      zz_rom_11[45] = 1'b1;
      zz_rom_11[46] = 1'b1;
      zz_rom_11[47] = 1'b1;
      zz_rom_11[48] = 1'b1;
      zz_rom_11[49] = 1'b1;
      zz_rom_11[50] = 1'b1;
      zz_rom_11[51] = 1'b1;
      zz_rom_11[52] = 1'b1;
      zz_rom_11[53] = 1'b1;
      zz_rom_11[54] = 1'b1;
      zz_rom_11[55] = 1'b1;
      zz_rom_11[56] = 1'b1;
      zz_rom_11[57] = 1'b1;
      zz_rom_11[58] = 1'b1;
      zz_rom_11[59] = 1'b1;
      zz_rom_11[60] = 1'b1;
      zz_rom_11[61] = 1'b1;
      zz_rom_11[62] = 1'b1;
      zz_rom_11[63] = 1'b1;
      zz_rom_11[64] = 1'b1;
      zz_rom_11[65] = 1'b1;
      zz_rom_11[66] = 1'b1;
      zz_rom_11[67] = 1'b1;
      zz_rom_11[68] = 1'b1;
      zz_rom_11[69] = 1'b1;
      zz_rom_11[70] = 1'b1;
      zz_rom_11[71] = 1'b1;
      zz_rom_11[72] = 1'b1;
      zz_rom_11[73] = 1'b1;
      zz_rom_11[74] = 1'b1;
      zz_rom_11[75] = 1'b1;
      zz_rom_11[76] = 1'b1;
      zz_rom_11[77] = 1'b1;
      zz_rom_11[78] = 1'b1;
      zz_rom_11[79] = 1'b1;
      zz_rom_11[80] = 1'b1;
      zz_rom_11[81] = 1'b1;
      zz_rom_11[82] = 1'b0;
      zz_rom_11[83] = 1'b0;
      zz_rom_11[84] = 1'b0;
      zz_rom_11[85] = 1'b0;
      zz_rom_11[86] = 1'b0;
      zz_rom_11[87] = 1'b0;
      zz_rom_11[88] = 1'b0;
      zz_rom_11[89] = 1'b0;
      zz_rom_11[90] = 1'b0;
      zz_rom_11[91] = 1'b0;
      zz_rom_11[92] = 1'b0;
      zz_rom_11[93] = 1'b0;
      zz_rom_11[94] = 1'b0;
      zz_rom_11[95] = 1'b0;
      zz_rom_11[96] = 1'b0;
      zz_rom_11[97] = 1'b0;
      zz_rom_11[98] = 1'b0;
      zz_rom_11[99] = 1'b0;
    end
  endfunction
  wire [99:0] _zz_12;
  function [99:0] zz_rom_12(input dummy);
    begin
      zz_rom_12[0] = 1'b0;
      zz_rom_12[1] = 1'b0;
      zz_rom_12[2] = 1'b0;
      zz_rom_12[3] = 1'b0;
      zz_rom_12[4] = 1'b0;
      zz_rom_12[5] = 1'b0;
      zz_rom_12[6] = 1'b0;
      zz_rom_12[7] = 1'b0;
      zz_rom_12[8] = 1'b0;
      zz_rom_12[9] = 1'b0;
      zz_rom_12[10] = 1'b0;
      zz_rom_12[11] = 1'b0;
      zz_rom_12[12] = 1'b0;
      zz_rom_12[13] = 1'b0;
      zz_rom_12[14] = 1'b0;
      zz_rom_12[15] = 1'b0;
      zz_rom_12[16] = 1'b0;
      zz_rom_12[17] = 1'b0;
      zz_rom_12[18] = 1'b1;
      zz_rom_12[19] = 1'b1;
      zz_rom_12[20] = 1'b1;
      zz_rom_12[21] = 1'b1;
      zz_rom_12[22] = 1'b1;
      zz_rom_12[23] = 1'b1;
      zz_rom_12[24] = 1'b1;
      zz_rom_12[25] = 1'b1;
      zz_rom_12[26] = 1'b1;
      zz_rom_12[27] = 1'b1;
      zz_rom_12[28] = 1'b1;
      zz_rom_12[29] = 1'b1;
      zz_rom_12[30] = 1'b1;
      zz_rom_12[31] = 1'b1;
      zz_rom_12[32] = 1'b1;
      zz_rom_12[33] = 1'b1;
      zz_rom_12[34] = 1'b1;
      zz_rom_12[35] = 1'b1;
      zz_rom_12[36] = 1'b1;
      zz_rom_12[37] = 1'b1;
      zz_rom_12[38] = 1'b1;
      zz_rom_12[39] = 1'b1;
      zz_rom_12[40] = 1'b1;
      zz_rom_12[41] = 1'b1;
      zz_rom_12[42] = 1'b1;
      zz_rom_12[43] = 1'b1;
      zz_rom_12[44] = 1'b1;
      zz_rom_12[45] = 1'b1;
      zz_rom_12[46] = 1'b1;
      zz_rom_12[47] = 1'b1;
      zz_rom_12[48] = 1'b1;
      zz_rom_12[49] = 1'b1;
      zz_rom_12[50] = 1'b1;
      zz_rom_12[51] = 1'b1;
      zz_rom_12[52] = 1'b1;
      zz_rom_12[53] = 1'b1;
      zz_rom_12[54] = 1'b1;
      zz_rom_12[55] = 1'b1;
      zz_rom_12[56] = 1'b1;
      zz_rom_12[57] = 1'b1;
      zz_rom_12[58] = 1'b1;
      zz_rom_12[59] = 1'b1;
      zz_rom_12[60] = 1'b1;
      zz_rom_12[61] = 1'b1;
      zz_rom_12[62] = 1'b1;
      zz_rom_12[63] = 1'b1;
      zz_rom_12[64] = 1'b1;
      zz_rom_12[65] = 1'b1;
      zz_rom_12[66] = 1'b1;
      zz_rom_12[67] = 1'b1;
      zz_rom_12[68] = 1'b1;
      zz_rom_12[69] = 1'b1;
      zz_rom_12[70] = 1'b1;
      zz_rom_12[71] = 1'b1;
      zz_rom_12[72] = 1'b1;
      zz_rom_12[73] = 1'b1;
      zz_rom_12[74] = 1'b1;
      zz_rom_12[75] = 1'b1;
      zz_rom_12[76] = 1'b1;
      zz_rom_12[77] = 1'b1;
      zz_rom_12[78] = 1'b1;
      zz_rom_12[79] = 1'b1;
      zz_rom_12[80] = 1'b1;
      zz_rom_12[81] = 1'b1;
      zz_rom_12[82] = 1'b1;
      zz_rom_12[83] = 1'b0;
      zz_rom_12[84] = 1'b0;
      zz_rom_12[85] = 1'b0;
      zz_rom_12[86] = 1'b0;
      zz_rom_12[87] = 1'b0;
      zz_rom_12[88] = 1'b0;
      zz_rom_12[89] = 1'b0;
      zz_rom_12[90] = 1'b0;
      zz_rom_12[91] = 1'b0;
      zz_rom_12[92] = 1'b0;
      zz_rom_12[93] = 1'b0;
      zz_rom_12[94] = 1'b0;
      zz_rom_12[95] = 1'b0;
      zz_rom_12[96] = 1'b0;
      zz_rom_12[97] = 1'b0;
      zz_rom_12[98] = 1'b0;
      zz_rom_12[99] = 1'b0;
    end
  endfunction
  wire [99:0] _zz_13;
  function [99:0] zz_rom_13(input dummy);
    begin
      zz_rom_13[0] = 1'b0;
      zz_rom_13[1] = 1'b0;
      zz_rom_13[2] = 1'b0;
      zz_rom_13[3] = 1'b0;
      zz_rom_13[4] = 1'b0;
      zz_rom_13[5] = 1'b0;
      zz_rom_13[6] = 1'b0;
      zz_rom_13[7] = 1'b0;
      zz_rom_13[8] = 1'b0;
      zz_rom_13[9] = 1'b0;
      zz_rom_13[10] = 1'b0;
      zz_rom_13[11] = 1'b0;
      zz_rom_13[12] = 1'b0;
      zz_rom_13[13] = 1'b0;
      zz_rom_13[14] = 1'b0;
      zz_rom_13[15] = 1'b0;
      zz_rom_13[16] = 1'b0;
      zz_rom_13[17] = 1'b1;
      zz_rom_13[18] = 1'b1;
      zz_rom_13[19] = 1'b1;
      zz_rom_13[20] = 1'b1;
      zz_rom_13[21] = 1'b1;
      zz_rom_13[22] = 1'b1;
      zz_rom_13[23] = 1'b1;
      zz_rom_13[24] = 1'b1;
      zz_rom_13[25] = 1'b1;
      zz_rom_13[26] = 1'b1;
      zz_rom_13[27] = 1'b1;
      zz_rom_13[28] = 1'b1;
      zz_rom_13[29] = 1'b1;
      zz_rom_13[30] = 1'b1;
      zz_rom_13[31] = 1'b1;
      zz_rom_13[32] = 1'b1;
      zz_rom_13[33] = 1'b1;
      zz_rom_13[34] = 1'b1;
      zz_rom_13[35] = 1'b1;
      zz_rom_13[36] = 1'b1;
      zz_rom_13[37] = 1'b1;
      zz_rom_13[38] = 1'b1;
      zz_rom_13[39] = 1'b1;
      zz_rom_13[40] = 1'b1;
      zz_rom_13[41] = 1'b1;
      zz_rom_13[42] = 1'b1;
      zz_rom_13[43] = 1'b1;
      zz_rom_13[44] = 1'b1;
      zz_rom_13[45] = 1'b1;
      zz_rom_13[46] = 1'b1;
      zz_rom_13[47] = 1'b1;
      zz_rom_13[48] = 1'b1;
      zz_rom_13[49] = 1'b1;
      zz_rom_13[50] = 1'b1;
      zz_rom_13[51] = 1'b1;
      zz_rom_13[52] = 1'b1;
      zz_rom_13[53] = 1'b1;
      zz_rom_13[54] = 1'b1;
      zz_rom_13[55] = 1'b1;
      zz_rom_13[56] = 1'b1;
      zz_rom_13[57] = 1'b1;
      zz_rom_13[58] = 1'b1;
      zz_rom_13[59] = 1'b1;
      zz_rom_13[60] = 1'b1;
      zz_rom_13[61] = 1'b1;
      zz_rom_13[62] = 1'b1;
      zz_rom_13[63] = 1'b1;
      zz_rom_13[64] = 1'b1;
      zz_rom_13[65] = 1'b1;
      zz_rom_13[66] = 1'b1;
      zz_rom_13[67] = 1'b1;
      zz_rom_13[68] = 1'b1;
      zz_rom_13[69] = 1'b1;
      zz_rom_13[70] = 1'b1;
      zz_rom_13[71] = 1'b1;
      zz_rom_13[72] = 1'b1;
      zz_rom_13[73] = 1'b1;
      zz_rom_13[74] = 1'b1;
      zz_rom_13[75] = 1'b1;
      zz_rom_13[76] = 1'b1;
      zz_rom_13[77] = 1'b1;
      zz_rom_13[78] = 1'b1;
      zz_rom_13[79] = 1'b1;
      zz_rom_13[80] = 1'b1;
      zz_rom_13[81] = 1'b1;
      zz_rom_13[82] = 1'b1;
      zz_rom_13[83] = 1'b1;
      zz_rom_13[84] = 1'b0;
      zz_rom_13[85] = 1'b0;
      zz_rom_13[86] = 1'b0;
      zz_rom_13[87] = 1'b0;
      zz_rom_13[88] = 1'b0;
      zz_rom_13[89] = 1'b0;
      zz_rom_13[90] = 1'b0;
      zz_rom_13[91] = 1'b0;
      zz_rom_13[92] = 1'b0;
      zz_rom_13[93] = 1'b0;
      zz_rom_13[94] = 1'b0;
      zz_rom_13[95] = 1'b0;
      zz_rom_13[96] = 1'b0;
      zz_rom_13[97] = 1'b0;
      zz_rom_13[98] = 1'b0;
      zz_rom_13[99] = 1'b0;
    end
  endfunction
  wire [99:0] _zz_14;
  function [99:0] zz_rom_14(input dummy);
    begin
      zz_rom_14[0] = 1'b0;
      zz_rom_14[1] = 1'b0;
      zz_rom_14[2] = 1'b0;
      zz_rom_14[3] = 1'b0;
      zz_rom_14[4] = 1'b0;
      zz_rom_14[5] = 1'b0;
      zz_rom_14[6] = 1'b0;
      zz_rom_14[7] = 1'b0;
      zz_rom_14[8] = 1'b0;
      zz_rom_14[9] = 1'b0;
      zz_rom_14[10] = 1'b0;
      zz_rom_14[11] = 1'b0;
      zz_rom_14[12] = 1'b0;
      zz_rom_14[13] = 1'b0;
      zz_rom_14[14] = 1'b0;
      zz_rom_14[15] = 1'b0;
      zz_rom_14[16] = 1'b1;
      zz_rom_14[17] = 1'b1;
      zz_rom_14[18] = 1'b1;
      zz_rom_14[19] = 1'b1;
      zz_rom_14[20] = 1'b1;
      zz_rom_14[21] = 1'b1;
      zz_rom_14[22] = 1'b1;
      zz_rom_14[23] = 1'b1;
      zz_rom_14[24] = 1'b1;
      zz_rom_14[25] = 1'b1;
      zz_rom_14[26] = 1'b1;
      zz_rom_14[27] = 1'b1;
      zz_rom_14[28] = 1'b1;
      zz_rom_14[29] = 1'b1;
      zz_rom_14[30] = 1'b1;
      zz_rom_14[31] = 1'b1;
      zz_rom_14[32] = 1'b1;
      zz_rom_14[33] = 1'b1;
      zz_rom_14[34] = 1'b1;
      zz_rom_14[35] = 1'b1;
      zz_rom_14[36] = 1'b1;
      zz_rom_14[37] = 1'b1;
      zz_rom_14[38] = 1'b1;
      zz_rom_14[39] = 1'b1;
      zz_rom_14[40] = 1'b1;
      zz_rom_14[41] = 1'b1;
      zz_rom_14[42] = 1'b1;
      zz_rom_14[43] = 1'b1;
      zz_rom_14[44] = 1'b1;
      zz_rom_14[45] = 1'b1;
      zz_rom_14[46] = 1'b1;
      zz_rom_14[47] = 1'b1;
      zz_rom_14[48] = 1'b1;
      zz_rom_14[49] = 1'b1;
      zz_rom_14[50] = 1'b1;
      zz_rom_14[51] = 1'b1;
      zz_rom_14[52] = 1'b1;
      zz_rom_14[53] = 1'b1;
      zz_rom_14[54] = 1'b1;
      zz_rom_14[55] = 1'b1;
      zz_rom_14[56] = 1'b1;
      zz_rom_14[57] = 1'b1;
      zz_rom_14[58] = 1'b1;
      zz_rom_14[59] = 1'b1;
      zz_rom_14[60] = 1'b1;
      zz_rom_14[61] = 1'b1;
      zz_rom_14[62] = 1'b1;
      zz_rom_14[63] = 1'b1;
      zz_rom_14[64] = 1'b1;
      zz_rom_14[65] = 1'b1;
      zz_rom_14[66] = 1'b1;
      zz_rom_14[67] = 1'b1;
      zz_rom_14[68] = 1'b1;
      zz_rom_14[69] = 1'b1;
      zz_rom_14[70] = 1'b1;
      zz_rom_14[71] = 1'b1;
      zz_rom_14[72] = 1'b1;
      zz_rom_14[73] = 1'b1;
      zz_rom_14[74] = 1'b1;
      zz_rom_14[75] = 1'b1;
      zz_rom_14[76] = 1'b1;
      zz_rom_14[77] = 1'b1;
      zz_rom_14[78] = 1'b1;
      zz_rom_14[79] = 1'b1;
      zz_rom_14[80] = 1'b1;
      zz_rom_14[81] = 1'b1;
      zz_rom_14[82] = 1'b1;
      zz_rom_14[83] = 1'b1;
      zz_rom_14[84] = 1'b1;
      zz_rom_14[85] = 1'b0;
      zz_rom_14[86] = 1'b0;
      zz_rom_14[87] = 1'b0;
      zz_rom_14[88] = 1'b0;
      zz_rom_14[89] = 1'b0;
      zz_rom_14[90] = 1'b0;
      zz_rom_14[91] = 1'b0;
      zz_rom_14[92] = 1'b0;
      zz_rom_14[93] = 1'b0;
      zz_rom_14[94] = 1'b0;
      zz_rom_14[95] = 1'b0;
      zz_rom_14[96] = 1'b0;
      zz_rom_14[97] = 1'b0;
      zz_rom_14[98] = 1'b0;
      zz_rom_14[99] = 1'b0;
    end
  endfunction
  wire [99:0] _zz_15;
  function [99:0] zz_rom_15(input dummy);
    begin
      zz_rom_15[0] = 1'b0;
      zz_rom_15[1] = 1'b0;
      zz_rom_15[2] = 1'b0;
      zz_rom_15[3] = 1'b0;
      zz_rom_15[4] = 1'b0;
      zz_rom_15[5] = 1'b0;
      zz_rom_15[6] = 1'b0;
      zz_rom_15[7] = 1'b0;
      zz_rom_15[8] = 1'b0;
      zz_rom_15[9] = 1'b0;
      zz_rom_15[10] = 1'b0;
      zz_rom_15[11] = 1'b0;
      zz_rom_15[12] = 1'b0;
      zz_rom_15[13] = 1'b0;
      zz_rom_15[14] = 1'b0;
      zz_rom_15[15] = 1'b1;
      zz_rom_15[16] = 1'b1;
      zz_rom_15[17] = 1'b1;
      zz_rom_15[18] = 1'b1;
      zz_rom_15[19] = 1'b1;
      zz_rom_15[20] = 1'b1;
      zz_rom_15[21] = 1'b1;
      zz_rom_15[22] = 1'b1;
      zz_rom_15[23] = 1'b1;
      zz_rom_15[24] = 1'b1;
      zz_rom_15[25] = 1'b1;
      zz_rom_15[26] = 1'b1;
      zz_rom_15[27] = 1'b1;
      zz_rom_15[28] = 1'b1;
      zz_rom_15[29] = 1'b1;
      zz_rom_15[30] = 1'b1;
      zz_rom_15[31] = 1'b1;
      zz_rom_15[32] = 1'b1;
      zz_rom_15[33] = 1'b1;
      zz_rom_15[34] = 1'b1;
      zz_rom_15[35] = 1'b1;
      zz_rom_15[36] = 1'b1;
      zz_rom_15[37] = 1'b1;
      zz_rom_15[38] = 1'b1;
      zz_rom_15[39] = 1'b1;
      zz_rom_15[40] = 1'b1;
      zz_rom_15[41] = 1'b1;
      zz_rom_15[42] = 1'b1;
      zz_rom_15[43] = 1'b1;
      zz_rom_15[44] = 1'b1;
      zz_rom_15[45] = 1'b1;
      zz_rom_15[46] = 1'b1;
      zz_rom_15[47] = 1'b1;
      zz_rom_15[48] = 1'b1;
      zz_rom_15[49] = 1'b1;
      zz_rom_15[50] = 1'b1;
      zz_rom_15[51] = 1'b1;
      zz_rom_15[52] = 1'b1;
      zz_rom_15[53] = 1'b1;
      zz_rom_15[54] = 1'b1;
      zz_rom_15[55] = 1'b1;
      zz_rom_15[56] = 1'b1;
      zz_rom_15[57] = 1'b1;
      zz_rom_15[58] = 1'b1;
      zz_rom_15[59] = 1'b1;
      zz_rom_15[60] = 1'b1;
      zz_rom_15[61] = 1'b1;
      zz_rom_15[62] = 1'b1;
      zz_rom_15[63] = 1'b1;
      zz_rom_15[64] = 1'b1;
      zz_rom_15[65] = 1'b1;
      zz_rom_15[66] = 1'b1;
      zz_rom_15[67] = 1'b1;
      zz_rom_15[68] = 1'b1;
      zz_rom_15[69] = 1'b1;
      zz_rom_15[70] = 1'b1;
      zz_rom_15[71] = 1'b1;
      zz_rom_15[72] = 1'b1;
      zz_rom_15[73] = 1'b1;
      zz_rom_15[74] = 1'b1;
      zz_rom_15[75] = 1'b1;
      zz_rom_15[76] = 1'b1;
      zz_rom_15[77] = 1'b1;
      zz_rom_15[78] = 1'b1;
      zz_rom_15[79] = 1'b1;
      zz_rom_15[80] = 1'b1;
      zz_rom_15[81] = 1'b1;
      zz_rom_15[82] = 1'b1;
      zz_rom_15[83] = 1'b1;
      zz_rom_15[84] = 1'b1;
      zz_rom_15[85] = 1'b1;
      zz_rom_15[86] = 1'b0;
      zz_rom_15[87] = 1'b0;
      zz_rom_15[88] = 1'b0;
      zz_rom_15[89] = 1'b0;
      zz_rom_15[90] = 1'b0;
      zz_rom_15[91] = 1'b0;
      zz_rom_15[92] = 1'b0;
      zz_rom_15[93] = 1'b0;
      zz_rom_15[94] = 1'b0;
      zz_rom_15[95] = 1'b0;
      zz_rom_15[96] = 1'b0;
      zz_rom_15[97] = 1'b0;
      zz_rom_15[98] = 1'b0;
      zz_rom_15[99] = 1'b0;
    end
  endfunction
  wire [99:0] _zz_16;
  function [99:0] zz_rom_16(input dummy);
    begin
      zz_rom_16[0] = 1'b0;
      zz_rom_16[1] = 1'b0;
      zz_rom_16[2] = 1'b0;
      zz_rom_16[3] = 1'b0;
      zz_rom_16[4] = 1'b0;
      zz_rom_16[5] = 1'b0;
      zz_rom_16[6] = 1'b0;
      zz_rom_16[7] = 1'b0;
      zz_rom_16[8] = 1'b0;
      zz_rom_16[9] = 1'b0;
      zz_rom_16[10] = 1'b0;
      zz_rom_16[11] = 1'b0;
      zz_rom_16[12] = 1'b0;
      zz_rom_16[13] = 1'b0;
      zz_rom_16[14] = 1'b1;
      zz_rom_16[15] = 1'b1;
      zz_rom_16[16] = 1'b1;
      zz_rom_16[17] = 1'b1;
      zz_rom_16[18] = 1'b1;
      zz_rom_16[19] = 1'b1;
      zz_rom_16[20] = 1'b1;
      zz_rom_16[21] = 1'b1;
      zz_rom_16[22] = 1'b1;
      zz_rom_16[23] = 1'b1;
      zz_rom_16[24] = 1'b1;
      zz_rom_16[25] = 1'b1;
      zz_rom_16[26] = 1'b1;
      zz_rom_16[27] = 1'b1;
      zz_rom_16[28] = 1'b1;
      zz_rom_16[29] = 1'b1;
      zz_rom_16[30] = 1'b1;
      zz_rom_16[31] = 1'b1;
      zz_rom_16[32] = 1'b1;
      zz_rom_16[33] = 1'b1;
      zz_rom_16[34] = 1'b1;
      zz_rom_16[35] = 1'b1;
      zz_rom_16[36] = 1'b1;
      zz_rom_16[37] = 1'b1;
      zz_rom_16[38] = 1'b1;
      zz_rom_16[39] = 1'b1;
      zz_rom_16[40] = 1'b1;
      zz_rom_16[41] = 1'b1;
      zz_rom_16[42] = 1'b1;
      zz_rom_16[43] = 1'b1;
      zz_rom_16[44] = 1'b1;
      zz_rom_16[45] = 1'b1;
      zz_rom_16[46] = 1'b1;
      zz_rom_16[47] = 1'b1;
      zz_rom_16[48] = 1'b1;
      zz_rom_16[49] = 1'b1;
      zz_rom_16[50] = 1'b1;
      zz_rom_16[51] = 1'b1;
      zz_rom_16[52] = 1'b1;
      zz_rom_16[53] = 1'b1;
      zz_rom_16[54] = 1'b1;
      zz_rom_16[55] = 1'b1;
      zz_rom_16[56] = 1'b1;
      zz_rom_16[57] = 1'b1;
      zz_rom_16[58] = 1'b1;
      zz_rom_16[59] = 1'b1;
      zz_rom_16[60] = 1'b1;
      zz_rom_16[61] = 1'b1;
      zz_rom_16[62] = 1'b1;
      zz_rom_16[63] = 1'b1;
      zz_rom_16[64] = 1'b1;
      zz_rom_16[65] = 1'b1;
      zz_rom_16[66] = 1'b1;
      zz_rom_16[67] = 1'b1;
      zz_rom_16[68] = 1'b1;
      zz_rom_16[69] = 1'b1;
      zz_rom_16[70] = 1'b1;
      zz_rom_16[71] = 1'b1;
      zz_rom_16[72] = 1'b1;
      zz_rom_16[73] = 1'b1;
      zz_rom_16[74] = 1'b1;
      zz_rom_16[75] = 1'b1;
      zz_rom_16[76] = 1'b1;
      zz_rom_16[77] = 1'b1;
      zz_rom_16[78] = 1'b1;
      zz_rom_16[79] = 1'b1;
      zz_rom_16[80] = 1'b1;
      zz_rom_16[81] = 1'b1;
      zz_rom_16[82] = 1'b1;
      zz_rom_16[83] = 1'b1;
      zz_rom_16[84] = 1'b1;
      zz_rom_16[85] = 1'b1;
      zz_rom_16[86] = 1'b1;
      zz_rom_16[87] = 1'b0;
      zz_rom_16[88] = 1'b0;
      zz_rom_16[89] = 1'b0;
      zz_rom_16[90] = 1'b0;
      zz_rom_16[91] = 1'b0;
      zz_rom_16[92] = 1'b0;
      zz_rom_16[93] = 1'b0;
      zz_rom_16[94] = 1'b0;
      zz_rom_16[95] = 1'b0;
      zz_rom_16[96] = 1'b0;
      zz_rom_16[97] = 1'b0;
      zz_rom_16[98] = 1'b0;
      zz_rom_16[99] = 1'b0;
    end
  endfunction
  wire [99:0] _zz_17;
  function [99:0] zz_rom_17(input dummy);
    begin
      zz_rom_17[0] = 1'b0;
      zz_rom_17[1] = 1'b0;
      zz_rom_17[2] = 1'b0;
      zz_rom_17[3] = 1'b0;
      zz_rom_17[4] = 1'b0;
      zz_rom_17[5] = 1'b0;
      zz_rom_17[6] = 1'b0;
      zz_rom_17[7] = 1'b0;
      zz_rom_17[8] = 1'b0;
      zz_rom_17[9] = 1'b0;
      zz_rom_17[10] = 1'b0;
      zz_rom_17[11] = 1'b0;
      zz_rom_17[12] = 1'b0;
      zz_rom_17[13] = 1'b1;
      zz_rom_17[14] = 1'b1;
      zz_rom_17[15] = 1'b1;
      zz_rom_17[16] = 1'b1;
      zz_rom_17[17] = 1'b1;
      zz_rom_17[18] = 1'b1;
      zz_rom_17[19] = 1'b1;
      zz_rom_17[20] = 1'b1;
      zz_rom_17[21] = 1'b1;
      zz_rom_17[22] = 1'b1;
      zz_rom_17[23] = 1'b1;
      zz_rom_17[24] = 1'b1;
      zz_rom_17[25] = 1'b1;
      zz_rom_17[26] = 1'b1;
      zz_rom_17[27] = 1'b1;
      zz_rom_17[28] = 1'b1;
      zz_rom_17[29] = 1'b1;
      zz_rom_17[30] = 1'b1;
      zz_rom_17[31] = 1'b1;
      zz_rom_17[32] = 1'b1;
      zz_rom_17[33] = 1'b1;
      zz_rom_17[34] = 1'b1;
      zz_rom_17[35] = 1'b1;
      zz_rom_17[36] = 1'b1;
      zz_rom_17[37] = 1'b1;
      zz_rom_17[38] = 1'b1;
      zz_rom_17[39] = 1'b1;
      zz_rom_17[40] = 1'b1;
      zz_rom_17[41] = 1'b1;
      zz_rom_17[42] = 1'b1;
      zz_rom_17[43] = 1'b1;
      zz_rom_17[44] = 1'b1;
      zz_rom_17[45] = 1'b1;
      zz_rom_17[46] = 1'b1;
      zz_rom_17[47] = 1'b1;
      zz_rom_17[48] = 1'b1;
      zz_rom_17[49] = 1'b1;
      zz_rom_17[50] = 1'b1;
      zz_rom_17[51] = 1'b1;
      zz_rom_17[52] = 1'b1;
      zz_rom_17[53] = 1'b1;
      zz_rom_17[54] = 1'b1;
      zz_rom_17[55] = 1'b1;
      zz_rom_17[56] = 1'b1;
      zz_rom_17[57] = 1'b1;
      zz_rom_17[58] = 1'b1;
      zz_rom_17[59] = 1'b1;
      zz_rom_17[60] = 1'b1;
      zz_rom_17[61] = 1'b1;
      zz_rom_17[62] = 1'b1;
      zz_rom_17[63] = 1'b1;
      zz_rom_17[64] = 1'b1;
      zz_rom_17[65] = 1'b1;
      zz_rom_17[66] = 1'b1;
      zz_rom_17[67] = 1'b1;
      zz_rom_17[68] = 1'b1;
      zz_rom_17[69] = 1'b1;
      zz_rom_17[70] = 1'b1;
      zz_rom_17[71] = 1'b1;
      zz_rom_17[72] = 1'b1;
      zz_rom_17[73] = 1'b1;
      zz_rom_17[74] = 1'b1;
      zz_rom_17[75] = 1'b1;
      zz_rom_17[76] = 1'b1;
      zz_rom_17[77] = 1'b1;
      zz_rom_17[78] = 1'b1;
      zz_rom_17[79] = 1'b1;
      zz_rom_17[80] = 1'b1;
      zz_rom_17[81] = 1'b1;
      zz_rom_17[82] = 1'b1;
      zz_rom_17[83] = 1'b1;
      zz_rom_17[84] = 1'b1;
      zz_rom_17[85] = 1'b1;
      zz_rom_17[86] = 1'b1;
      zz_rom_17[87] = 1'b1;
      zz_rom_17[88] = 1'b0;
      zz_rom_17[89] = 1'b0;
      zz_rom_17[90] = 1'b0;
      zz_rom_17[91] = 1'b0;
      zz_rom_17[92] = 1'b0;
      zz_rom_17[93] = 1'b0;
      zz_rom_17[94] = 1'b0;
      zz_rom_17[95] = 1'b0;
      zz_rom_17[96] = 1'b0;
      zz_rom_17[97] = 1'b0;
      zz_rom_17[98] = 1'b0;
      zz_rom_17[99] = 1'b0;
    end
  endfunction
  wire [99:0] _zz_18;
  function [99:0] zz_rom_18(input dummy);
    begin
      zz_rom_18[0] = 1'b0;
      zz_rom_18[1] = 1'b0;
      zz_rom_18[2] = 1'b0;
      zz_rom_18[3] = 1'b0;
      zz_rom_18[4] = 1'b0;
      zz_rom_18[5] = 1'b0;
      zz_rom_18[6] = 1'b0;
      zz_rom_18[7] = 1'b0;
      zz_rom_18[8] = 1'b0;
      zz_rom_18[9] = 1'b0;
      zz_rom_18[10] = 1'b0;
      zz_rom_18[11] = 1'b0;
      zz_rom_18[12] = 1'b1;
      zz_rom_18[13] = 1'b1;
      zz_rom_18[14] = 1'b1;
      zz_rom_18[15] = 1'b1;
      zz_rom_18[16] = 1'b1;
      zz_rom_18[17] = 1'b1;
      zz_rom_18[18] = 1'b1;
      zz_rom_18[19] = 1'b1;
      zz_rom_18[20] = 1'b1;
      zz_rom_18[21] = 1'b1;
      zz_rom_18[22] = 1'b1;
      zz_rom_18[23] = 1'b1;
      zz_rom_18[24] = 1'b1;
      zz_rom_18[25] = 1'b1;
      zz_rom_18[26] = 1'b1;
      zz_rom_18[27] = 1'b1;
      zz_rom_18[28] = 1'b1;
      zz_rom_18[29] = 1'b1;
      zz_rom_18[30] = 1'b1;
      zz_rom_18[31] = 1'b1;
      zz_rom_18[32] = 1'b1;
      zz_rom_18[33] = 1'b1;
      zz_rom_18[34] = 1'b1;
      zz_rom_18[35] = 1'b1;
      zz_rom_18[36] = 1'b1;
      zz_rom_18[37] = 1'b1;
      zz_rom_18[38] = 1'b1;
      zz_rom_18[39] = 1'b1;
      zz_rom_18[40] = 1'b1;
      zz_rom_18[41] = 1'b1;
      zz_rom_18[42] = 1'b1;
      zz_rom_18[43] = 1'b1;
      zz_rom_18[44] = 1'b1;
      zz_rom_18[45] = 1'b1;
      zz_rom_18[46] = 1'b1;
      zz_rom_18[47] = 1'b1;
      zz_rom_18[48] = 1'b1;
      zz_rom_18[49] = 1'b1;
      zz_rom_18[50] = 1'b1;
      zz_rom_18[51] = 1'b1;
      zz_rom_18[52] = 1'b1;
      zz_rom_18[53] = 1'b1;
      zz_rom_18[54] = 1'b1;
      zz_rom_18[55] = 1'b1;
      zz_rom_18[56] = 1'b1;
      zz_rom_18[57] = 1'b1;
      zz_rom_18[58] = 1'b1;
      zz_rom_18[59] = 1'b1;
      zz_rom_18[60] = 1'b1;
      zz_rom_18[61] = 1'b1;
      zz_rom_18[62] = 1'b1;
      zz_rom_18[63] = 1'b1;
      zz_rom_18[64] = 1'b1;
      zz_rom_18[65] = 1'b1;
      zz_rom_18[66] = 1'b1;
      zz_rom_18[67] = 1'b1;
      zz_rom_18[68] = 1'b1;
      zz_rom_18[69] = 1'b1;
      zz_rom_18[70] = 1'b1;
      zz_rom_18[71] = 1'b1;
      zz_rom_18[72] = 1'b1;
      zz_rom_18[73] = 1'b1;
      zz_rom_18[74] = 1'b1;
      zz_rom_18[75] = 1'b1;
      zz_rom_18[76] = 1'b1;
      zz_rom_18[77] = 1'b1;
      zz_rom_18[78] = 1'b1;
      zz_rom_18[79] = 1'b1;
      zz_rom_18[80] = 1'b1;
      zz_rom_18[81] = 1'b1;
      zz_rom_18[82] = 1'b1;
      zz_rom_18[83] = 1'b1;
      zz_rom_18[84] = 1'b1;
      zz_rom_18[85] = 1'b1;
      zz_rom_18[86] = 1'b1;
      zz_rom_18[87] = 1'b1;
      zz_rom_18[88] = 1'b1;
      zz_rom_18[89] = 1'b0;
      zz_rom_18[90] = 1'b0;
      zz_rom_18[91] = 1'b0;
      zz_rom_18[92] = 1'b0;
      zz_rom_18[93] = 1'b0;
      zz_rom_18[94] = 1'b0;
      zz_rom_18[95] = 1'b0;
      zz_rom_18[96] = 1'b0;
      zz_rom_18[97] = 1'b0;
      zz_rom_18[98] = 1'b0;
      zz_rom_18[99] = 1'b0;
    end
  endfunction
  wire [99:0] _zz_19;
  function [99:0] zz_rom_19(input dummy);
    begin
      zz_rom_19[0] = 1'b0;
      zz_rom_19[1] = 1'b0;
      zz_rom_19[2] = 1'b0;
      zz_rom_19[3] = 1'b0;
      zz_rom_19[4] = 1'b0;
      zz_rom_19[5] = 1'b0;
      zz_rom_19[6] = 1'b0;
      zz_rom_19[7] = 1'b0;
      zz_rom_19[8] = 1'b0;
      zz_rom_19[9] = 1'b0;
      zz_rom_19[10] = 1'b0;
      zz_rom_19[11] = 1'b1;
      zz_rom_19[12] = 1'b1;
      zz_rom_19[13] = 1'b1;
      zz_rom_19[14] = 1'b1;
      zz_rom_19[15] = 1'b1;
      zz_rom_19[16] = 1'b1;
      zz_rom_19[17] = 1'b1;
      zz_rom_19[18] = 1'b1;
      zz_rom_19[19] = 1'b1;
      zz_rom_19[20] = 1'b1;
      zz_rom_19[21] = 1'b1;
      zz_rom_19[22] = 1'b1;
      zz_rom_19[23] = 1'b1;
      zz_rom_19[24] = 1'b1;
      zz_rom_19[25] = 1'b1;
      zz_rom_19[26] = 1'b1;
      zz_rom_19[27] = 1'b1;
      zz_rom_19[28] = 1'b1;
      zz_rom_19[29] = 1'b1;
      zz_rom_19[30] = 1'b1;
      zz_rom_19[31] = 1'b1;
      zz_rom_19[32] = 1'b1;
      zz_rom_19[33] = 1'b1;
      zz_rom_19[34] = 1'b1;
      zz_rom_19[35] = 1'b1;
      zz_rom_19[36] = 1'b1;
      zz_rom_19[37] = 1'b1;
      zz_rom_19[38] = 1'b1;
      zz_rom_19[39] = 1'b1;
      zz_rom_19[40] = 1'b1;
      zz_rom_19[41] = 1'b1;
      zz_rom_19[42] = 1'b1;
      zz_rom_19[43] = 1'b1;
      zz_rom_19[44] = 1'b1;
      zz_rom_19[45] = 1'b1;
      zz_rom_19[46] = 1'b1;
      zz_rom_19[47] = 1'b1;
      zz_rom_19[48] = 1'b1;
      zz_rom_19[49] = 1'b1;
      zz_rom_19[50] = 1'b1;
      zz_rom_19[51] = 1'b1;
      zz_rom_19[52] = 1'b1;
      zz_rom_19[53] = 1'b1;
      zz_rom_19[54] = 1'b1;
      zz_rom_19[55] = 1'b1;
      zz_rom_19[56] = 1'b1;
      zz_rom_19[57] = 1'b1;
      zz_rom_19[58] = 1'b1;
      zz_rom_19[59] = 1'b1;
      zz_rom_19[60] = 1'b1;
      zz_rom_19[61] = 1'b1;
      zz_rom_19[62] = 1'b1;
      zz_rom_19[63] = 1'b1;
      zz_rom_19[64] = 1'b1;
      zz_rom_19[65] = 1'b1;
      zz_rom_19[66] = 1'b1;
      zz_rom_19[67] = 1'b1;
      zz_rom_19[68] = 1'b1;
      zz_rom_19[69] = 1'b1;
      zz_rom_19[70] = 1'b1;
      zz_rom_19[71] = 1'b1;
      zz_rom_19[72] = 1'b1;
      zz_rom_19[73] = 1'b1;
      zz_rom_19[74] = 1'b1;
      zz_rom_19[75] = 1'b1;
      zz_rom_19[76] = 1'b1;
      zz_rom_19[77] = 1'b1;
      zz_rom_19[78] = 1'b1;
      zz_rom_19[79] = 1'b1;
      zz_rom_19[80] = 1'b1;
      zz_rom_19[81] = 1'b1;
      zz_rom_19[82] = 1'b1;
      zz_rom_19[83] = 1'b1;
      zz_rom_19[84] = 1'b1;
      zz_rom_19[85] = 1'b1;
      zz_rom_19[86] = 1'b1;
      zz_rom_19[87] = 1'b1;
      zz_rom_19[88] = 1'b1;
      zz_rom_19[89] = 1'b1;
      zz_rom_19[90] = 1'b0;
      zz_rom_19[91] = 1'b0;
      zz_rom_19[92] = 1'b0;
      zz_rom_19[93] = 1'b0;
      zz_rom_19[94] = 1'b0;
      zz_rom_19[95] = 1'b0;
      zz_rom_19[96] = 1'b0;
      zz_rom_19[97] = 1'b0;
      zz_rom_19[98] = 1'b0;
      zz_rom_19[99] = 1'b0;
    end
  endfunction
  wire [99:0] _zz_20;
  function [99:0] zz_rom_20(input dummy);
    begin
      zz_rom_20[0] = 1'b0;
      zz_rom_20[1] = 1'b0;
      zz_rom_20[2] = 1'b0;
      zz_rom_20[3] = 1'b0;
      zz_rom_20[4] = 1'b0;
      zz_rom_20[5] = 1'b0;
      zz_rom_20[6] = 1'b0;
      zz_rom_20[7] = 1'b0;
      zz_rom_20[8] = 1'b0;
      zz_rom_20[9] = 1'b0;
      zz_rom_20[10] = 1'b1;
      zz_rom_20[11] = 1'b1;
      zz_rom_20[12] = 1'b1;
      zz_rom_20[13] = 1'b1;
      zz_rom_20[14] = 1'b1;
      zz_rom_20[15] = 1'b1;
      zz_rom_20[16] = 1'b1;
      zz_rom_20[17] = 1'b1;
      zz_rom_20[18] = 1'b1;
      zz_rom_20[19] = 1'b1;
      zz_rom_20[20] = 1'b1;
      zz_rom_20[21] = 1'b1;
      zz_rom_20[22] = 1'b1;
      zz_rom_20[23] = 1'b1;
      zz_rom_20[24] = 1'b1;
      zz_rom_20[25] = 1'b1;
      zz_rom_20[26] = 1'b1;
      zz_rom_20[27] = 1'b1;
      zz_rom_20[28] = 1'b1;
      zz_rom_20[29] = 1'b1;
      zz_rom_20[30] = 1'b1;
      zz_rom_20[31] = 1'b1;
      zz_rom_20[32] = 1'b1;
      zz_rom_20[33] = 1'b1;
      zz_rom_20[34] = 1'b1;
      zz_rom_20[35] = 1'b1;
      zz_rom_20[36] = 1'b1;
      zz_rom_20[37] = 1'b1;
      zz_rom_20[38] = 1'b1;
      zz_rom_20[39] = 1'b1;
      zz_rom_20[40] = 1'b1;
      zz_rom_20[41] = 1'b1;
      zz_rom_20[42] = 1'b1;
      zz_rom_20[43] = 1'b1;
      zz_rom_20[44] = 1'b1;
      zz_rom_20[45] = 1'b1;
      zz_rom_20[46] = 1'b1;
      zz_rom_20[47] = 1'b1;
      zz_rom_20[48] = 1'b1;
      zz_rom_20[49] = 1'b1;
      zz_rom_20[50] = 1'b1;
      zz_rom_20[51] = 1'b1;
      zz_rom_20[52] = 1'b1;
      zz_rom_20[53] = 1'b1;
      zz_rom_20[54] = 1'b1;
      zz_rom_20[55] = 1'b1;
      zz_rom_20[56] = 1'b1;
      zz_rom_20[57] = 1'b1;
      zz_rom_20[58] = 1'b1;
      zz_rom_20[59] = 1'b1;
      zz_rom_20[60] = 1'b1;
      zz_rom_20[61] = 1'b1;
      zz_rom_20[62] = 1'b1;
      zz_rom_20[63] = 1'b1;
      zz_rom_20[64] = 1'b1;
      zz_rom_20[65] = 1'b1;
      zz_rom_20[66] = 1'b1;
      zz_rom_20[67] = 1'b1;
      zz_rom_20[68] = 1'b1;
      zz_rom_20[69] = 1'b1;
      zz_rom_20[70] = 1'b1;
      zz_rom_20[71] = 1'b1;
      zz_rom_20[72] = 1'b1;
      zz_rom_20[73] = 1'b1;
      zz_rom_20[74] = 1'b1;
      zz_rom_20[75] = 1'b1;
      zz_rom_20[76] = 1'b1;
      zz_rom_20[77] = 1'b1;
      zz_rom_20[78] = 1'b1;
      zz_rom_20[79] = 1'b1;
      zz_rom_20[80] = 1'b1;
      zz_rom_20[81] = 1'b1;
      zz_rom_20[82] = 1'b1;
      zz_rom_20[83] = 1'b1;
      zz_rom_20[84] = 1'b1;
      zz_rom_20[85] = 1'b1;
      zz_rom_20[86] = 1'b1;
      zz_rom_20[87] = 1'b1;
      zz_rom_20[88] = 1'b1;
      zz_rom_20[89] = 1'b1;
      zz_rom_20[90] = 1'b1;
      zz_rom_20[91] = 1'b0;
      zz_rom_20[92] = 1'b0;
      zz_rom_20[93] = 1'b0;
      zz_rom_20[94] = 1'b0;
      zz_rom_20[95] = 1'b0;
      zz_rom_20[96] = 1'b0;
      zz_rom_20[97] = 1'b0;
      zz_rom_20[98] = 1'b0;
      zz_rom_20[99] = 1'b0;
    end
  endfunction
  wire [99:0] _zz_21;
  function [99:0] zz_rom_21(input dummy);
    begin
      zz_rom_21[0] = 1'b0;
      zz_rom_21[1] = 1'b0;
      zz_rom_21[2] = 1'b0;
      zz_rom_21[3] = 1'b0;
      zz_rom_21[4] = 1'b0;
      zz_rom_21[5] = 1'b0;
      zz_rom_21[6] = 1'b0;
      zz_rom_21[7] = 1'b0;
      zz_rom_21[8] = 1'b0;
      zz_rom_21[9] = 1'b0;
      zz_rom_21[10] = 1'b1;
      zz_rom_21[11] = 1'b1;
      zz_rom_21[12] = 1'b1;
      zz_rom_21[13] = 1'b1;
      zz_rom_21[14] = 1'b1;
      zz_rom_21[15] = 1'b1;
      zz_rom_21[16] = 1'b1;
      zz_rom_21[17] = 1'b1;
      zz_rom_21[18] = 1'b1;
      zz_rom_21[19] = 1'b1;
      zz_rom_21[20] = 1'b1;
      zz_rom_21[21] = 1'b1;
      zz_rom_21[22] = 1'b1;
      zz_rom_21[23] = 1'b1;
      zz_rom_21[24] = 1'b1;
      zz_rom_21[25] = 1'b1;
      zz_rom_21[26] = 1'b1;
      zz_rom_21[27] = 1'b1;
      zz_rom_21[28] = 1'b1;
      zz_rom_21[29] = 1'b1;
      zz_rom_21[30] = 1'b1;
      zz_rom_21[31] = 1'b1;
      zz_rom_21[32] = 1'b1;
      zz_rom_21[33] = 1'b1;
      zz_rom_21[34] = 1'b1;
      zz_rom_21[35] = 1'b1;
      zz_rom_21[36] = 1'b1;
      zz_rom_21[37] = 1'b1;
      zz_rom_21[38] = 1'b1;
      zz_rom_21[39] = 1'b1;
      zz_rom_21[40] = 1'b1;
      zz_rom_21[41] = 1'b1;
      zz_rom_21[42] = 1'b1;
      zz_rom_21[43] = 1'b1;
      zz_rom_21[44] = 1'b1;
      zz_rom_21[45] = 1'b1;
      zz_rom_21[46] = 1'b1;
      zz_rom_21[47] = 1'b1;
      zz_rom_21[48] = 1'b1;
      zz_rom_21[49] = 1'b1;
      zz_rom_21[50] = 1'b1;
      zz_rom_21[51] = 1'b1;
      zz_rom_21[52] = 1'b1;
      zz_rom_21[53] = 1'b1;
      zz_rom_21[54] = 1'b1;
      zz_rom_21[55] = 1'b1;
      zz_rom_21[56] = 1'b1;
      zz_rom_21[57] = 1'b1;
      zz_rom_21[58] = 1'b1;
      zz_rom_21[59] = 1'b1;
      zz_rom_21[60] = 1'b1;
      zz_rom_21[61] = 1'b1;
      zz_rom_21[62] = 1'b1;
      zz_rom_21[63] = 1'b1;
      zz_rom_21[64] = 1'b1;
      zz_rom_21[65] = 1'b1;
      zz_rom_21[66] = 1'b1;
      zz_rom_21[67] = 1'b1;
      zz_rom_21[68] = 1'b1;
      zz_rom_21[69] = 1'b1;
      zz_rom_21[70] = 1'b1;
      zz_rom_21[71] = 1'b1;
      zz_rom_21[72] = 1'b1;
      zz_rom_21[73] = 1'b1;
      zz_rom_21[74] = 1'b1;
      zz_rom_21[75] = 1'b1;
      zz_rom_21[76] = 1'b1;
      zz_rom_21[77] = 1'b1;
      zz_rom_21[78] = 1'b1;
      zz_rom_21[79] = 1'b1;
      zz_rom_21[80] = 1'b1;
      zz_rom_21[81] = 1'b1;
      zz_rom_21[82] = 1'b1;
      zz_rom_21[83] = 1'b1;
      zz_rom_21[84] = 1'b1;
      zz_rom_21[85] = 1'b1;
      zz_rom_21[86] = 1'b1;
      zz_rom_21[87] = 1'b1;
      zz_rom_21[88] = 1'b1;
      zz_rom_21[89] = 1'b1;
      zz_rom_21[90] = 1'b1;
      zz_rom_21[91] = 1'b0;
      zz_rom_21[92] = 1'b0;
      zz_rom_21[93] = 1'b0;
      zz_rom_21[94] = 1'b0;
      zz_rom_21[95] = 1'b0;
      zz_rom_21[96] = 1'b0;
      zz_rom_21[97] = 1'b0;
      zz_rom_21[98] = 1'b0;
      zz_rom_21[99] = 1'b0;
    end
  endfunction
  wire [99:0] _zz_22;
  function [99:0] zz_rom_22(input dummy);
    begin
      zz_rom_22[0] = 1'b0;
      zz_rom_22[1] = 1'b0;
      zz_rom_22[2] = 1'b0;
      zz_rom_22[3] = 1'b0;
      zz_rom_22[4] = 1'b0;
      zz_rom_22[5] = 1'b0;
      zz_rom_22[6] = 1'b0;
      zz_rom_22[7] = 1'b0;
      zz_rom_22[8] = 1'b0;
      zz_rom_22[9] = 1'b1;
      zz_rom_22[10] = 1'b1;
      zz_rom_22[11] = 1'b1;
      zz_rom_22[12] = 1'b1;
      zz_rom_22[13] = 1'b1;
      zz_rom_22[14] = 1'b1;
      zz_rom_22[15] = 1'b1;
      zz_rom_22[16] = 1'b1;
      zz_rom_22[17] = 1'b1;
      zz_rom_22[18] = 1'b1;
      zz_rom_22[19] = 1'b1;
      zz_rom_22[20] = 1'b1;
      zz_rom_22[21] = 1'b1;
      zz_rom_22[22] = 1'b1;
      zz_rom_22[23] = 1'b1;
      zz_rom_22[24] = 1'b1;
      zz_rom_22[25] = 1'b1;
      zz_rom_22[26] = 1'b1;
      zz_rom_22[27] = 1'b1;
      zz_rom_22[28] = 1'b1;
      zz_rom_22[29] = 1'b1;
      zz_rom_22[30] = 1'b1;
      zz_rom_22[31] = 1'b1;
      zz_rom_22[32] = 1'b1;
      zz_rom_22[33] = 1'b1;
      zz_rom_22[34] = 1'b1;
      zz_rom_22[35] = 1'b1;
      zz_rom_22[36] = 1'b1;
      zz_rom_22[37] = 1'b1;
      zz_rom_22[38] = 1'b1;
      zz_rom_22[39] = 1'b1;
      zz_rom_22[40] = 1'b1;
      zz_rom_22[41] = 1'b1;
      zz_rom_22[42] = 1'b1;
      zz_rom_22[43] = 1'b1;
      zz_rom_22[44] = 1'b1;
      zz_rom_22[45] = 1'b1;
      zz_rom_22[46] = 1'b1;
      zz_rom_22[47] = 1'b1;
      zz_rom_22[48] = 1'b1;
      zz_rom_22[49] = 1'b1;
      zz_rom_22[50] = 1'b1;
      zz_rom_22[51] = 1'b1;
      zz_rom_22[52] = 1'b1;
      zz_rom_22[53] = 1'b1;
      zz_rom_22[54] = 1'b1;
      zz_rom_22[55] = 1'b1;
      zz_rom_22[56] = 1'b1;
      zz_rom_22[57] = 1'b1;
      zz_rom_22[58] = 1'b1;
      zz_rom_22[59] = 1'b1;
      zz_rom_22[60] = 1'b1;
      zz_rom_22[61] = 1'b1;
      zz_rom_22[62] = 1'b1;
      zz_rom_22[63] = 1'b1;
      zz_rom_22[64] = 1'b1;
      zz_rom_22[65] = 1'b1;
      zz_rom_22[66] = 1'b1;
      zz_rom_22[67] = 1'b1;
      zz_rom_22[68] = 1'b1;
      zz_rom_22[69] = 1'b1;
      zz_rom_22[70] = 1'b1;
      zz_rom_22[71] = 1'b1;
      zz_rom_22[72] = 1'b1;
      zz_rom_22[73] = 1'b1;
      zz_rom_22[74] = 1'b1;
      zz_rom_22[75] = 1'b1;
      zz_rom_22[76] = 1'b1;
      zz_rom_22[77] = 1'b1;
      zz_rom_22[78] = 1'b1;
      zz_rom_22[79] = 1'b1;
      zz_rom_22[80] = 1'b1;
      zz_rom_22[81] = 1'b1;
      zz_rom_22[82] = 1'b1;
      zz_rom_22[83] = 1'b1;
      zz_rom_22[84] = 1'b1;
      zz_rom_22[85] = 1'b1;
      zz_rom_22[86] = 1'b1;
      zz_rom_22[87] = 1'b1;
      zz_rom_22[88] = 1'b1;
      zz_rom_22[89] = 1'b1;
      zz_rom_22[90] = 1'b1;
      zz_rom_22[91] = 1'b1;
      zz_rom_22[92] = 1'b0;
      zz_rom_22[93] = 1'b0;
      zz_rom_22[94] = 1'b0;
      zz_rom_22[95] = 1'b0;
      zz_rom_22[96] = 1'b0;
      zz_rom_22[97] = 1'b0;
      zz_rom_22[98] = 1'b0;
      zz_rom_22[99] = 1'b0;
    end
  endfunction
  wire [99:0] _zz_23;
  function [99:0] zz_rom_23(input dummy);
    begin
      zz_rom_23[0] = 1'b0;
      zz_rom_23[1] = 1'b0;
      zz_rom_23[2] = 1'b0;
      zz_rom_23[3] = 1'b0;
      zz_rom_23[4] = 1'b0;
      zz_rom_23[5] = 1'b0;
      zz_rom_23[6] = 1'b0;
      zz_rom_23[7] = 1'b0;
      zz_rom_23[8] = 1'b1;
      zz_rom_23[9] = 1'b1;
      zz_rom_23[10] = 1'b1;
      zz_rom_23[11] = 1'b1;
      zz_rom_23[12] = 1'b1;
      zz_rom_23[13] = 1'b1;
      zz_rom_23[14] = 1'b1;
      zz_rom_23[15] = 1'b1;
      zz_rom_23[16] = 1'b1;
      zz_rom_23[17] = 1'b1;
      zz_rom_23[18] = 1'b1;
      zz_rom_23[19] = 1'b1;
      zz_rom_23[20] = 1'b1;
      zz_rom_23[21] = 1'b1;
      zz_rom_23[22] = 1'b1;
      zz_rom_23[23] = 1'b1;
      zz_rom_23[24] = 1'b1;
      zz_rom_23[25] = 1'b1;
      zz_rom_23[26] = 1'b1;
      zz_rom_23[27] = 1'b1;
      zz_rom_23[28] = 1'b1;
      zz_rom_23[29] = 1'b1;
      zz_rom_23[30] = 1'b1;
      zz_rom_23[31] = 1'b1;
      zz_rom_23[32] = 1'b1;
      zz_rom_23[33] = 1'b1;
      zz_rom_23[34] = 1'b1;
      zz_rom_23[35] = 1'b1;
      zz_rom_23[36] = 1'b1;
      zz_rom_23[37] = 1'b1;
      zz_rom_23[38] = 1'b1;
      zz_rom_23[39] = 1'b1;
      zz_rom_23[40] = 1'b1;
      zz_rom_23[41] = 1'b1;
      zz_rom_23[42] = 1'b1;
      zz_rom_23[43] = 1'b1;
      zz_rom_23[44] = 1'b1;
      zz_rom_23[45] = 1'b1;
      zz_rom_23[46] = 1'b1;
      zz_rom_23[47] = 1'b1;
      zz_rom_23[48] = 1'b1;
      zz_rom_23[49] = 1'b1;
      zz_rom_23[50] = 1'b1;
      zz_rom_23[51] = 1'b1;
      zz_rom_23[52] = 1'b1;
      zz_rom_23[53] = 1'b1;
      zz_rom_23[54] = 1'b1;
      zz_rom_23[55] = 1'b1;
      zz_rom_23[56] = 1'b1;
      zz_rom_23[57] = 1'b1;
      zz_rom_23[58] = 1'b1;
      zz_rom_23[59] = 1'b1;
      zz_rom_23[60] = 1'b1;
      zz_rom_23[61] = 1'b1;
      zz_rom_23[62] = 1'b1;
      zz_rom_23[63] = 1'b1;
      zz_rom_23[64] = 1'b1;
      zz_rom_23[65] = 1'b1;
      zz_rom_23[66] = 1'b1;
      zz_rom_23[67] = 1'b1;
      zz_rom_23[68] = 1'b1;
      zz_rom_23[69] = 1'b1;
      zz_rom_23[70] = 1'b1;
      zz_rom_23[71] = 1'b1;
      zz_rom_23[72] = 1'b1;
      zz_rom_23[73] = 1'b1;
      zz_rom_23[74] = 1'b1;
      zz_rom_23[75] = 1'b1;
      zz_rom_23[76] = 1'b1;
      zz_rom_23[77] = 1'b1;
      zz_rom_23[78] = 1'b1;
      zz_rom_23[79] = 1'b1;
      zz_rom_23[80] = 1'b1;
      zz_rom_23[81] = 1'b1;
      zz_rom_23[82] = 1'b1;
      zz_rom_23[83] = 1'b1;
      zz_rom_23[84] = 1'b1;
      zz_rom_23[85] = 1'b1;
      zz_rom_23[86] = 1'b1;
      zz_rom_23[87] = 1'b1;
      zz_rom_23[88] = 1'b1;
      zz_rom_23[89] = 1'b1;
      zz_rom_23[90] = 1'b1;
      zz_rom_23[91] = 1'b1;
      zz_rom_23[92] = 1'b1;
      zz_rom_23[93] = 1'b0;
      zz_rom_23[94] = 1'b0;
      zz_rom_23[95] = 1'b0;
      zz_rom_23[96] = 1'b0;
      zz_rom_23[97] = 1'b0;
      zz_rom_23[98] = 1'b0;
      zz_rom_23[99] = 1'b0;
    end
  endfunction
  wire [99:0] _zz_24;
  function [99:0] zz_rom_24(input dummy);
    begin
      zz_rom_24[0] = 1'b0;
      zz_rom_24[1] = 1'b0;
      zz_rom_24[2] = 1'b0;
      zz_rom_24[3] = 1'b0;
      zz_rom_24[4] = 1'b0;
      zz_rom_24[5] = 1'b0;
      zz_rom_24[6] = 1'b0;
      zz_rom_24[7] = 1'b0;
      zz_rom_24[8] = 1'b1;
      zz_rom_24[9] = 1'b1;
      zz_rom_24[10] = 1'b1;
      zz_rom_24[11] = 1'b1;
      zz_rom_24[12] = 1'b1;
      zz_rom_24[13] = 1'b1;
      zz_rom_24[14] = 1'b1;
      zz_rom_24[15] = 1'b1;
      zz_rom_24[16] = 1'b1;
      zz_rom_24[17] = 1'b1;
      zz_rom_24[18] = 1'b1;
      zz_rom_24[19] = 1'b1;
      zz_rom_24[20] = 1'b1;
      zz_rom_24[21] = 1'b1;
      zz_rom_24[22] = 1'b1;
      zz_rom_24[23] = 1'b1;
      zz_rom_24[24] = 1'b1;
      zz_rom_24[25] = 1'b1;
      zz_rom_24[26] = 1'b1;
      zz_rom_24[27] = 1'b1;
      zz_rom_24[28] = 1'b1;
      zz_rom_24[29] = 1'b1;
      zz_rom_24[30] = 1'b1;
      zz_rom_24[31] = 1'b1;
      zz_rom_24[32] = 1'b1;
      zz_rom_24[33] = 1'b1;
      zz_rom_24[34] = 1'b1;
      zz_rom_24[35] = 1'b1;
      zz_rom_24[36] = 1'b1;
      zz_rom_24[37] = 1'b1;
      zz_rom_24[38] = 1'b1;
      zz_rom_24[39] = 1'b1;
      zz_rom_24[40] = 1'b1;
      zz_rom_24[41] = 1'b1;
      zz_rom_24[42] = 1'b1;
      zz_rom_24[43] = 1'b1;
      zz_rom_24[44] = 1'b1;
      zz_rom_24[45] = 1'b1;
      zz_rom_24[46] = 1'b1;
      zz_rom_24[47] = 1'b1;
      zz_rom_24[48] = 1'b1;
      zz_rom_24[49] = 1'b1;
      zz_rom_24[50] = 1'b1;
      zz_rom_24[51] = 1'b1;
      zz_rom_24[52] = 1'b1;
      zz_rom_24[53] = 1'b1;
      zz_rom_24[54] = 1'b1;
      zz_rom_24[55] = 1'b1;
      zz_rom_24[56] = 1'b1;
      zz_rom_24[57] = 1'b1;
      zz_rom_24[58] = 1'b1;
      zz_rom_24[59] = 1'b1;
      zz_rom_24[60] = 1'b1;
      zz_rom_24[61] = 1'b1;
      zz_rom_24[62] = 1'b1;
      zz_rom_24[63] = 1'b1;
      zz_rom_24[64] = 1'b1;
      zz_rom_24[65] = 1'b1;
      zz_rom_24[66] = 1'b1;
      zz_rom_24[67] = 1'b1;
      zz_rom_24[68] = 1'b1;
      zz_rom_24[69] = 1'b1;
      zz_rom_24[70] = 1'b1;
      zz_rom_24[71] = 1'b1;
      zz_rom_24[72] = 1'b1;
      zz_rom_24[73] = 1'b1;
      zz_rom_24[74] = 1'b1;
      zz_rom_24[75] = 1'b1;
      zz_rom_24[76] = 1'b1;
      zz_rom_24[77] = 1'b1;
      zz_rom_24[78] = 1'b1;
      zz_rom_24[79] = 1'b1;
      zz_rom_24[80] = 1'b1;
      zz_rom_24[81] = 1'b1;
      zz_rom_24[82] = 1'b1;
      zz_rom_24[83] = 1'b1;
      zz_rom_24[84] = 1'b1;
      zz_rom_24[85] = 1'b1;
      zz_rom_24[86] = 1'b1;
      zz_rom_24[87] = 1'b1;
      zz_rom_24[88] = 1'b1;
      zz_rom_24[89] = 1'b1;
      zz_rom_24[90] = 1'b1;
      zz_rom_24[91] = 1'b1;
      zz_rom_24[92] = 1'b1;
      zz_rom_24[93] = 1'b0;
      zz_rom_24[94] = 1'b0;
      zz_rom_24[95] = 1'b0;
      zz_rom_24[96] = 1'b0;
      zz_rom_24[97] = 1'b0;
      zz_rom_24[98] = 1'b0;
      zz_rom_24[99] = 1'b0;
    end
  endfunction
  wire [99:0] _zz_25;
  function [99:0] zz_rom_25(input dummy);
    begin
      zz_rom_25[0] = 1'b0;
      zz_rom_25[1] = 1'b0;
      zz_rom_25[2] = 1'b0;
      zz_rom_25[3] = 1'b0;
      zz_rom_25[4] = 1'b0;
      zz_rom_25[5] = 1'b0;
      zz_rom_25[6] = 1'b0;
      zz_rom_25[7] = 1'b1;
      zz_rom_25[8] = 1'b1;
      zz_rom_25[9] = 1'b1;
      zz_rom_25[10] = 1'b1;
      zz_rom_25[11] = 1'b1;
      zz_rom_25[12] = 1'b1;
      zz_rom_25[13] = 1'b1;
      zz_rom_25[14] = 1'b1;
      zz_rom_25[15] = 1'b1;
      zz_rom_25[16] = 1'b1;
      zz_rom_25[17] = 1'b1;
      zz_rom_25[18] = 1'b1;
      zz_rom_25[19] = 1'b1;
      zz_rom_25[20] = 1'b1;
      zz_rom_25[21] = 1'b1;
      zz_rom_25[22] = 1'b1;
      zz_rom_25[23] = 1'b1;
      zz_rom_25[24] = 1'b1;
      zz_rom_25[25] = 1'b1;
      zz_rom_25[26] = 1'b1;
      zz_rom_25[27] = 1'b1;
      zz_rom_25[28] = 1'b1;
      zz_rom_25[29] = 1'b1;
      zz_rom_25[30] = 1'b1;
      zz_rom_25[31] = 1'b1;
      zz_rom_25[32] = 1'b1;
      zz_rom_25[33] = 1'b1;
      zz_rom_25[34] = 1'b1;
      zz_rom_25[35] = 1'b1;
      zz_rom_25[36] = 1'b1;
      zz_rom_25[37] = 1'b1;
      zz_rom_25[38] = 1'b1;
      zz_rom_25[39] = 1'b1;
      zz_rom_25[40] = 1'b1;
      zz_rom_25[41] = 1'b1;
      zz_rom_25[42] = 1'b1;
      zz_rom_25[43] = 1'b1;
      zz_rom_25[44] = 1'b1;
      zz_rom_25[45] = 1'b1;
      zz_rom_25[46] = 1'b1;
      zz_rom_25[47] = 1'b1;
      zz_rom_25[48] = 1'b1;
      zz_rom_25[49] = 1'b1;
      zz_rom_25[50] = 1'b1;
      zz_rom_25[51] = 1'b1;
      zz_rom_25[52] = 1'b1;
      zz_rom_25[53] = 1'b1;
      zz_rom_25[54] = 1'b1;
      zz_rom_25[55] = 1'b1;
      zz_rom_25[56] = 1'b1;
      zz_rom_25[57] = 1'b1;
      zz_rom_25[58] = 1'b1;
      zz_rom_25[59] = 1'b1;
      zz_rom_25[60] = 1'b1;
      zz_rom_25[61] = 1'b1;
      zz_rom_25[62] = 1'b1;
      zz_rom_25[63] = 1'b1;
      zz_rom_25[64] = 1'b1;
      zz_rom_25[65] = 1'b1;
      zz_rom_25[66] = 1'b1;
      zz_rom_25[67] = 1'b1;
      zz_rom_25[68] = 1'b1;
      zz_rom_25[69] = 1'b1;
      zz_rom_25[70] = 1'b1;
      zz_rom_25[71] = 1'b1;
      zz_rom_25[72] = 1'b1;
      zz_rom_25[73] = 1'b1;
      zz_rom_25[74] = 1'b1;
      zz_rom_25[75] = 1'b1;
      zz_rom_25[76] = 1'b1;
      zz_rom_25[77] = 1'b1;
      zz_rom_25[78] = 1'b1;
      zz_rom_25[79] = 1'b1;
      zz_rom_25[80] = 1'b1;
      zz_rom_25[81] = 1'b1;
      zz_rom_25[82] = 1'b1;
      zz_rom_25[83] = 1'b1;
      zz_rom_25[84] = 1'b1;
      zz_rom_25[85] = 1'b1;
      zz_rom_25[86] = 1'b1;
      zz_rom_25[87] = 1'b1;
      zz_rom_25[88] = 1'b1;
      zz_rom_25[89] = 1'b1;
      zz_rom_25[90] = 1'b1;
      zz_rom_25[91] = 1'b1;
      zz_rom_25[92] = 1'b1;
      zz_rom_25[93] = 1'b1;
      zz_rom_25[94] = 1'b0;
      zz_rom_25[95] = 1'b0;
      zz_rom_25[96] = 1'b0;
      zz_rom_25[97] = 1'b0;
      zz_rom_25[98] = 1'b0;
      zz_rom_25[99] = 1'b0;
    end
  endfunction
  wire [99:0] _zz_26;
  function [99:0] zz_rom_26(input dummy);
    begin
      zz_rom_26[0] = 1'b0;
      zz_rom_26[1] = 1'b0;
      zz_rom_26[2] = 1'b0;
      zz_rom_26[3] = 1'b0;
      zz_rom_26[4] = 1'b0;
      zz_rom_26[5] = 1'b0;
      zz_rom_26[6] = 1'b0;
      zz_rom_26[7] = 1'b1;
      zz_rom_26[8] = 1'b1;
      zz_rom_26[9] = 1'b1;
      zz_rom_26[10] = 1'b1;
      zz_rom_26[11] = 1'b1;
      zz_rom_26[12] = 1'b1;
      zz_rom_26[13] = 1'b1;
      zz_rom_26[14] = 1'b1;
      zz_rom_26[15] = 1'b1;
      zz_rom_26[16] = 1'b1;
      zz_rom_26[17] = 1'b1;
      zz_rom_26[18] = 1'b1;
      zz_rom_26[19] = 1'b1;
      zz_rom_26[20] = 1'b1;
      zz_rom_26[21] = 1'b1;
      zz_rom_26[22] = 1'b1;
      zz_rom_26[23] = 1'b1;
      zz_rom_26[24] = 1'b1;
      zz_rom_26[25] = 1'b1;
      zz_rom_26[26] = 1'b1;
      zz_rom_26[27] = 1'b1;
      zz_rom_26[28] = 1'b1;
      zz_rom_26[29] = 1'b1;
      zz_rom_26[30] = 1'b1;
      zz_rom_26[31] = 1'b1;
      zz_rom_26[32] = 1'b1;
      zz_rom_26[33] = 1'b1;
      zz_rom_26[34] = 1'b1;
      zz_rom_26[35] = 1'b1;
      zz_rom_26[36] = 1'b1;
      zz_rom_26[37] = 1'b1;
      zz_rom_26[38] = 1'b1;
      zz_rom_26[39] = 1'b1;
      zz_rom_26[40] = 1'b1;
      zz_rom_26[41] = 1'b1;
      zz_rom_26[42] = 1'b1;
      zz_rom_26[43] = 1'b1;
      zz_rom_26[44] = 1'b1;
      zz_rom_26[45] = 1'b1;
      zz_rom_26[46] = 1'b1;
      zz_rom_26[47] = 1'b1;
      zz_rom_26[48] = 1'b1;
      zz_rom_26[49] = 1'b1;
      zz_rom_26[50] = 1'b1;
      zz_rom_26[51] = 1'b1;
      zz_rom_26[52] = 1'b1;
      zz_rom_26[53] = 1'b1;
      zz_rom_26[54] = 1'b1;
      zz_rom_26[55] = 1'b1;
      zz_rom_26[56] = 1'b1;
      zz_rom_26[57] = 1'b1;
      zz_rom_26[58] = 1'b1;
      zz_rom_26[59] = 1'b1;
      zz_rom_26[60] = 1'b1;
      zz_rom_26[61] = 1'b1;
      zz_rom_26[62] = 1'b1;
      zz_rom_26[63] = 1'b1;
      zz_rom_26[64] = 1'b1;
      zz_rom_26[65] = 1'b1;
      zz_rom_26[66] = 1'b1;
      zz_rom_26[67] = 1'b1;
      zz_rom_26[68] = 1'b1;
      zz_rom_26[69] = 1'b1;
      zz_rom_26[70] = 1'b1;
      zz_rom_26[71] = 1'b1;
      zz_rom_26[72] = 1'b1;
      zz_rom_26[73] = 1'b1;
      zz_rom_26[74] = 1'b1;
      zz_rom_26[75] = 1'b1;
      zz_rom_26[76] = 1'b1;
      zz_rom_26[77] = 1'b1;
      zz_rom_26[78] = 1'b1;
      zz_rom_26[79] = 1'b1;
      zz_rom_26[80] = 1'b1;
      zz_rom_26[81] = 1'b1;
      zz_rom_26[82] = 1'b1;
      zz_rom_26[83] = 1'b1;
      zz_rom_26[84] = 1'b1;
      zz_rom_26[85] = 1'b1;
      zz_rom_26[86] = 1'b1;
      zz_rom_26[87] = 1'b1;
      zz_rom_26[88] = 1'b1;
      zz_rom_26[89] = 1'b1;
      zz_rom_26[90] = 1'b1;
      zz_rom_26[91] = 1'b1;
      zz_rom_26[92] = 1'b1;
      zz_rom_26[93] = 1'b1;
      zz_rom_26[94] = 1'b0;
      zz_rom_26[95] = 1'b0;
      zz_rom_26[96] = 1'b0;
      zz_rom_26[97] = 1'b0;
      zz_rom_26[98] = 1'b0;
      zz_rom_26[99] = 1'b0;
    end
  endfunction
  wire [99:0] _zz_27;
  function [99:0] zz_rom_27(input dummy);
    begin
      zz_rom_27[0] = 1'b0;
      zz_rom_27[1] = 1'b0;
      zz_rom_27[2] = 1'b0;
      zz_rom_27[3] = 1'b0;
      zz_rom_27[4] = 1'b0;
      zz_rom_27[5] = 1'b0;
      zz_rom_27[6] = 1'b1;
      zz_rom_27[7] = 1'b1;
      zz_rom_27[8] = 1'b1;
      zz_rom_27[9] = 1'b1;
      zz_rom_27[10] = 1'b1;
      zz_rom_27[11] = 1'b1;
      zz_rom_27[12] = 1'b1;
      zz_rom_27[13] = 1'b1;
      zz_rom_27[14] = 1'b1;
      zz_rom_27[15] = 1'b1;
      zz_rom_27[16] = 1'b1;
      zz_rom_27[17] = 1'b1;
      zz_rom_27[18] = 1'b1;
      zz_rom_27[19] = 1'b1;
      zz_rom_27[20] = 1'b1;
      zz_rom_27[21] = 1'b1;
      zz_rom_27[22] = 1'b1;
      zz_rom_27[23] = 1'b1;
      zz_rom_27[24] = 1'b1;
      zz_rom_27[25] = 1'b1;
      zz_rom_27[26] = 1'b1;
      zz_rom_27[27] = 1'b1;
      zz_rom_27[28] = 1'b1;
      zz_rom_27[29] = 1'b1;
      zz_rom_27[30] = 1'b1;
      zz_rom_27[31] = 1'b1;
      zz_rom_27[32] = 1'b1;
      zz_rom_27[33] = 1'b1;
      zz_rom_27[34] = 1'b1;
      zz_rom_27[35] = 1'b1;
      zz_rom_27[36] = 1'b1;
      zz_rom_27[37] = 1'b1;
      zz_rom_27[38] = 1'b1;
      zz_rom_27[39] = 1'b1;
      zz_rom_27[40] = 1'b1;
      zz_rom_27[41] = 1'b1;
      zz_rom_27[42] = 1'b1;
      zz_rom_27[43] = 1'b1;
      zz_rom_27[44] = 1'b1;
      zz_rom_27[45] = 1'b1;
      zz_rom_27[46] = 1'b1;
      zz_rom_27[47] = 1'b1;
      zz_rom_27[48] = 1'b1;
      zz_rom_27[49] = 1'b1;
      zz_rom_27[50] = 1'b1;
      zz_rom_27[51] = 1'b1;
      zz_rom_27[52] = 1'b1;
      zz_rom_27[53] = 1'b1;
      zz_rom_27[54] = 1'b1;
      zz_rom_27[55] = 1'b1;
      zz_rom_27[56] = 1'b1;
      zz_rom_27[57] = 1'b1;
      zz_rom_27[58] = 1'b1;
      zz_rom_27[59] = 1'b1;
      zz_rom_27[60] = 1'b1;
      zz_rom_27[61] = 1'b1;
      zz_rom_27[62] = 1'b1;
      zz_rom_27[63] = 1'b1;
      zz_rom_27[64] = 1'b1;
      zz_rom_27[65] = 1'b1;
      zz_rom_27[66] = 1'b1;
      zz_rom_27[67] = 1'b1;
      zz_rom_27[68] = 1'b1;
      zz_rom_27[69] = 1'b1;
      zz_rom_27[70] = 1'b1;
      zz_rom_27[71] = 1'b1;
      zz_rom_27[72] = 1'b1;
      zz_rom_27[73] = 1'b1;
      zz_rom_27[74] = 1'b1;
      zz_rom_27[75] = 1'b1;
      zz_rom_27[76] = 1'b1;
      zz_rom_27[77] = 1'b1;
      zz_rom_27[78] = 1'b1;
      zz_rom_27[79] = 1'b1;
      zz_rom_27[80] = 1'b1;
      zz_rom_27[81] = 1'b1;
      zz_rom_27[82] = 1'b1;
      zz_rom_27[83] = 1'b1;
      zz_rom_27[84] = 1'b1;
      zz_rom_27[85] = 1'b1;
      zz_rom_27[86] = 1'b1;
      zz_rom_27[87] = 1'b1;
      zz_rom_27[88] = 1'b1;
      zz_rom_27[89] = 1'b1;
      zz_rom_27[90] = 1'b1;
      zz_rom_27[91] = 1'b1;
      zz_rom_27[92] = 1'b1;
      zz_rom_27[93] = 1'b1;
      zz_rom_27[94] = 1'b1;
      zz_rom_27[95] = 1'b0;
      zz_rom_27[96] = 1'b0;
      zz_rom_27[97] = 1'b0;
      zz_rom_27[98] = 1'b0;
      zz_rom_27[99] = 1'b0;
    end
  endfunction
  wire [99:0] _zz_28;
  function [99:0] zz_rom_28(input dummy);
    begin
      zz_rom_28[0] = 1'b0;
      zz_rom_28[1] = 1'b0;
      zz_rom_28[2] = 1'b0;
      zz_rom_28[3] = 1'b0;
      zz_rom_28[4] = 1'b0;
      zz_rom_28[5] = 1'b0;
      zz_rom_28[6] = 1'b1;
      zz_rom_28[7] = 1'b1;
      zz_rom_28[8] = 1'b1;
      zz_rom_28[9] = 1'b1;
      zz_rom_28[10] = 1'b1;
      zz_rom_28[11] = 1'b1;
      zz_rom_28[12] = 1'b1;
      zz_rom_28[13] = 1'b1;
      zz_rom_28[14] = 1'b1;
      zz_rom_28[15] = 1'b1;
      zz_rom_28[16] = 1'b1;
      zz_rom_28[17] = 1'b1;
      zz_rom_28[18] = 1'b1;
      zz_rom_28[19] = 1'b1;
      zz_rom_28[20] = 1'b1;
      zz_rom_28[21] = 1'b1;
      zz_rom_28[22] = 1'b1;
      zz_rom_28[23] = 1'b1;
      zz_rom_28[24] = 1'b1;
      zz_rom_28[25] = 1'b1;
      zz_rom_28[26] = 1'b1;
      zz_rom_28[27] = 1'b1;
      zz_rom_28[28] = 1'b1;
      zz_rom_28[29] = 1'b1;
      zz_rom_28[30] = 1'b1;
      zz_rom_28[31] = 1'b1;
      zz_rom_28[32] = 1'b1;
      zz_rom_28[33] = 1'b1;
      zz_rom_28[34] = 1'b1;
      zz_rom_28[35] = 1'b1;
      zz_rom_28[36] = 1'b1;
      zz_rom_28[37] = 1'b1;
      zz_rom_28[38] = 1'b1;
      zz_rom_28[39] = 1'b1;
      zz_rom_28[40] = 1'b1;
      zz_rom_28[41] = 1'b1;
      zz_rom_28[42] = 1'b1;
      zz_rom_28[43] = 1'b1;
      zz_rom_28[44] = 1'b1;
      zz_rom_28[45] = 1'b1;
      zz_rom_28[46] = 1'b1;
      zz_rom_28[47] = 1'b1;
      zz_rom_28[48] = 1'b1;
      zz_rom_28[49] = 1'b1;
      zz_rom_28[50] = 1'b1;
      zz_rom_28[51] = 1'b1;
      zz_rom_28[52] = 1'b1;
      zz_rom_28[53] = 1'b1;
      zz_rom_28[54] = 1'b1;
      zz_rom_28[55] = 1'b1;
      zz_rom_28[56] = 1'b1;
      zz_rom_28[57] = 1'b1;
      zz_rom_28[58] = 1'b1;
      zz_rom_28[59] = 1'b1;
      zz_rom_28[60] = 1'b1;
      zz_rom_28[61] = 1'b1;
      zz_rom_28[62] = 1'b1;
      zz_rom_28[63] = 1'b1;
      zz_rom_28[64] = 1'b1;
      zz_rom_28[65] = 1'b1;
      zz_rom_28[66] = 1'b1;
      zz_rom_28[67] = 1'b1;
      zz_rom_28[68] = 1'b1;
      zz_rom_28[69] = 1'b1;
      zz_rom_28[70] = 1'b1;
      zz_rom_28[71] = 1'b1;
      zz_rom_28[72] = 1'b1;
      zz_rom_28[73] = 1'b1;
      zz_rom_28[74] = 1'b1;
      zz_rom_28[75] = 1'b1;
      zz_rom_28[76] = 1'b1;
      zz_rom_28[77] = 1'b1;
      zz_rom_28[78] = 1'b1;
      zz_rom_28[79] = 1'b1;
      zz_rom_28[80] = 1'b1;
      zz_rom_28[81] = 1'b1;
      zz_rom_28[82] = 1'b1;
      zz_rom_28[83] = 1'b1;
      zz_rom_28[84] = 1'b1;
      zz_rom_28[85] = 1'b1;
      zz_rom_28[86] = 1'b1;
      zz_rom_28[87] = 1'b1;
      zz_rom_28[88] = 1'b1;
      zz_rom_28[89] = 1'b1;
      zz_rom_28[90] = 1'b1;
      zz_rom_28[91] = 1'b1;
      zz_rom_28[92] = 1'b1;
      zz_rom_28[93] = 1'b1;
      zz_rom_28[94] = 1'b1;
      zz_rom_28[95] = 1'b0;
      zz_rom_28[96] = 1'b0;
      zz_rom_28[97] = 1'b0;
      zz_rom_28[98] = 1'b0;
      zz_rom_28[99] = 1'b0;
    end
  endfunction
  wire [99:0] _zz_29;
  function [99:0] zz_rom_29(input dummy);
    begin
      zz_rom_29[0] = 1'b0;
      zz_rom_29[1] = 1'b0;
      zz_rom_29[2] = 1'b0;
      zz_rom_29[3] = 1'b0;
      zz_rom_29[4] = 1'b0;
      zz_rom_29[5] = 1'b1;
      zz_rom_29[6] = 1'b1;
      zz_rom_29[7] = 1'b1;
      zz_rom_29[8] = 1'b1;
      zz_rom_29[9] = 1'b1;
      zz_rom_29[10] = 1'b1;
      zz_rom_29[11] = 1'b1;
      zz_rom_29[12] = 1'b1;
      zz_rom_29[13] = 1'b1;
      zz_rom_29[14] = 1'b1;
      zz_rom_29[15] = 1'b1;
      zz_rom_29[16] = 1'b1;
      zz_rom_29[17] = 1'b1;
      zz_rom_29[18] = 1'b1;
      zz_rom_29[19] = 1'b1;
      zz_rom_29[20] = 1'b1;
      zz_rom_29[21] = 1'b1;
      zz_rom_29[22] = 1'b1;
      zz_rom_29[23] = 1'b1;
      zz_rom_29[24] = 1'b1;
      zz_rom_29[25] = 1'b1;
      zz_rom_29[26] = 1'b1;
      zz_rom_29[27] = 1'b1;
      zz_rom_29[28] = 1'b1;
      zz_rom_29[29] = 1'b1;
      zz_rom_29[30] = 1'b1;
      zz_rom_29[31] = 1'b1;
      zz_rom_29[32] = 1'b1;
      zz_rom_29[33] = 1'b1;
      zz_rom_29[34] = 1'b1;
      zz_rom_29[35] = 1'b1;
      zz_rom_29[36] = 1'b1;
      zz_rom_29[37] = 1'b1;
      zz_rom_29[38] = 1'b1;
      zz_rom_29[39] = 1'b1;
      zz_rom_29[40] = 1'b1;
      zz_rom_29[41] = 1'b1;
      zz_rom_29[42] = 1'b1;
      zz_rom_29[43] = 1'b1;
      zz_rom_29[44] = 1'b1;
      zz_rom_29[45] = 1'b1;
      zz_rom_29[46] = 1'b1;
      zz_rom_29[47] = 1'b1;
      zz_rom_29[48] = 1'b1;
      zz_rom_29[49] = 1'b1;
      zz_rom_29[50] = 1'b1;
      zz_rom_29[51] = 1'b1;
      zz_rom_29[52] = 1'b1;
      zz_rom_29[53] = 1'b1;
      zz_rom_29[54] = 1'b1;
      zz_rom_29[55] = 1'b1;
      zz_rom_29[56] = 1'b1;
      zz_rom_29[57] = 1'b1;
      zz_rom_29[58] = 1'b1;
      zz_rom_29[59] = 1'b1;
      zz_rom_29[60] = 1'b1;
      zz_rom_29[61] = 1'b1;
      zz_rom_29[62] = 1'b1;
      zz_rom_29[63] = 1'b1;
      zz_rom_29[64] = 1'b1;
      zz_rom_29[65] = 1'b1;
      zz_rom_29[66] = 1'b1;
      zz_rom_29[67] = 1'b1;
      zz_rom_29[68] = 1'b1;
      zz_rom_29[69] = 1'b1;
      zz_rom_29[70] = 1'b1;
      zz_rom_29[71] = 1'b1;
      zz_rom_29[72] = 1'b1;
      zz_rom_29[73] = 1'b1;
      zz_rom_29[74] = 1'b1;
      zz_rom_29[75] = 1'b1;
      zz_rom_29[76] = 1'b1;
      zz_rom_29[77] = 1'b1;
      zz_rom_29[78] = 1'b1;
      zz_rom_29[79] = 1'b1;
      zz_rom_29[80] = 1'b1;
      zz_rom_29[81] = 1'b1;
      zz_rom_29[82] = 1'b1;
      zz_rom_29[83] = 1'b1;
      zz_rom_29[84] = 1'b1;
      zz_rom_29[85] = 1'b1;
      zz_rom_29[86] = 1'b1;
      zz_rom_29[87] = 1'b1;
      zz_rom_29[88] = 1'b1;
      zz_rom_29[89] = 1'b1;
      zz_rom_29[90] = 1'b1;
      zz_rom_29[91] = 1'b1;
      zz_rom_29[92] = 1'b1;
      zz_rom_29[93] = 1'b1;
      zz_rom_29[94] = 1'b1;
      zz_rom_29[95] = 1'b1;
      zz_rom_29[96] = 1'b0;
      zz_rom_29[97] = 1'b0;
      zz_rom_29[98] = 1'b0;
      zz_rom_29[99] = 1'b0;
    end
  endfunction
  wire [99:0] _zz_30;
  function [99:0] zz_rom_30(input dummy);
    begin
      zz_rom_30[0] = 1'b0;
      zz_rom_30[1] = 1'b0;
      zz_rom_30[2] = 1'b0;
      zz_rom_30[3] = 1'b0;
      zz_rom_30[4] = 1'b0;
      zz_rom_30[5] = 1'b1;
      zz_rom_30[6] = 1'b1;
      zz_rom_30[7] = 1'b1;
      zz_rom_30[8] = 1'b1;
      zz_rom_30[9] = 1'b1;
      zz_rom_30[10] = 1'b1;
      zz_rom_30[11] = 1'b1;
      zz_rom_30[12] = 1'b1;
      zz_rom_30[13] = 1'b1;
      zz_rom_30[14] = 1'b1;
      zz_rom_30[15] = 1'b1;
      zz_rom_30[16] = 1'b1;
      zz_rom_30[17] = 1'b1;
      zz_rom_30[18] = 1'b1;
      zz_rom_30[19] = 1'b1;
      zz_rom_30[20] = 1'b1;
      zz_rom_30[21] = 1'b1;
      zz_rom_30[22] = 1'b1;
      zz_rom_30[23] = 1'b1;
      zz_rom_30[24] = 1'b1;
      zz_rom_30[25] = 1'b1;
      zz_rom_30[26] = 1'b1;
      zz_rom_30[27] = 1'b1;
      zz_rom_30[28] = 1'b1;
      zz_rom_30[29] = 1'b1;
      zz_rom_30[30] = 1'b1;
      zz_rom_30[31] = 1'b1;
      zz_rom_30[32] = 1'b1;
      zz_rom_30[33] = 1'b1;
      zz_rom_30[34] = 1'b1;
      zz_rom_30[35] = 1'b1;
      zz_rom_30[36] = 1'b1;
      zz_rom_30[37] = 1'b1;
      zz_rom_30[38] = 1'b1;
      zz_rom_30[39] = 1'b1;
      zz_rom_30[40] = 1'b1;
      zz_rom_30[41] = 1'b1;
      zz_rom_30[42] = 1'b1;
      zz_rom_30[43] = 1'b1;
      zz_rom_30[44] = 1'b1;
      zz_rom_30[45] = 1'b1;
      zz_rom_30[46] = 1'b1;
      zz_rom_30[47] = 1'b1;
      zz_rom_30[48] = 1'b1;
      zz_rom_30[49] = 1'b1;
      zz_rom_30[50] = 1'b1;
      zz_rom_30[51] = 1'b1;
      zz_rom_30[52] = 1'b1;
      zz_rom_30[53] = 1'b1;
      zz_rom_30[54] = 1'b1;
      zz_rom_30[55] = 1'b1;
      zz_rom_30[56] = 1'b1;
      zz_rom_30[57] = 1'b1;
      zz_rom_30[58] = 1'b1;
      zz_rom_30[59] = 1'b1;
      zz_rom_30[60] = 1'b1;
      zz_rom_30[61] = 1'b1;
      zz_rom_30[62] = 1'b1;
      zz_rom_30[63] = 1'b1;
      zz_rom_30[64] = 1'b1;
      zz_rom_30[65] = 1'b1;
      zz_rom_30[66] = 1'b1;
      zz_rom_30[67] = 1'b1;
      zz_rom_30[68] = 1'b1;
      zz_rom_30[69] = 1'b1;
      zz_rom_30[70] = 1'b1;
      zz_rom_30[71] = 1'b1;
      zz_rom_30[72] = 1'b1;
      zz_rom_30[73] = 1'b1;
      zz_rom_30[74] = 1'b1;
      zz_rom_30[75] = 1'b1;
      zz_rom_30[76] = 1'b1;
      zz_rom_30[77] = 1'b1;
      zz_rom_30[78] = 1'b1;
      zz_rom_30[79] = 1'b1;
      zz_rom_30[80] = 1'b1;
      zz_rom_30[81] = 1'b1;
      zz_rom_30[82] = 1'b1;
      zz_rom_30[83] = 1'b1;
      zz_rom_30[84] = 1'b1;
      zz_rom_30[85] = 1'b1;
      zz_rom_30[86] = 1'b1;
      zz_rom_30[87] = 1'b1;
      zz_rom_30[88] = 1'b1;
      zz_rom_30[89] = 1'b1;
      zz_rom_30[90] = 1'b1;
      zz_rom_30[91] = 1'b1;
      zz_rom_30[92] = 1'b1;
      zz_rom_30[93] = 1'b1;
      zz_rom_30[94] = 1'b1;
      zz_rom_30[95] = 1'b1;
      zz_rom_30[96] = 1'b0;
      zz_rom_30[97] = 1'b0;
      zz_rom_30[98] = 1'b0;
      zz_rom_30[99] = 1'b0;
    end
  endfunction
  wire [99:0] _zz_31;
  function [99:0] zz_rom_31(input dummy);
    begin
      zz_rom_31[0] = 1'b0;
      zz_rom_31[1] = 1'b0;
      zz_rom_31[2] = 1'b0;
      zz_rom_31[3] = 1'b0;
      zz_rom_31[4] = 1'b1;
      zz_rom_31[5] = 1'b1;
      zz_rom_31[6] = 1'b1;
      zz_rom_31[7] = 1'b1;
      zz_rom_31[8] = 1'b1;
      zz_rom_31[9] = 1'b1;
      zz_rom_31[10] = 1'b1;
      zz_rom_31[11] = 1'b1;
      zz_rom_31[12] = 1'b1;
      zz_rom_31[13] = 1'b1;
      zz_rom_31[14] = 1'b1;
      zz_rom_31[15] = 1'b1;
      zz_rom_31[16] = 1'b1;
      zz_rom_31[17] = 1'b1;
      zz_rom_31[18] = 1'b1;
      zz_rom_31[19] = 1'b1;
      zz_rom_31[20] = 1'b1;
      zz_rom_31[21] = 1'b1;
      zz_rom_31[22] = 1'b1;
      zz_rom_31[23] = 1'b1;
      zz_rom_31[24] = 1'b1;
      zz_rom_31[25] = 1'b1;
      zz_rom_31[26] = 1'b1;
      zz_rom_31[27] = 1'b1;
      zz_rom_31[28] = 1'b1;
      zz_rom_31[29] = 1'b1;
      zz_rom_31[30] = 1'b1;
      zz_rom_31[31] = 1'b1;
      zz_rom_31[32] = 1'b1;
      zz_rom_31[33] = 1'b1;
      zz_rom_31[34] = 1'b1;
      zz_rom_31[35] = 1'b1;
      zz_rom_31[36] = 1'b1;
      zz_rom_31[37] = 1'b1;
      zz_rom_31[38] = 1'b1;
      zz_rom_31[39] = 1'b1;
      zz_rom_31[40] = 1'b1;
      zz_rom_31[41] = 1'b1;
      zz_rom_31[42] = 1'b1;
      zz_rom_31[43] = 1'b1;
      zz_rom_31[44] = 1'b1;
      zz_rom_31[45] = 1'b1;
      zz_rom_31[46] = 1'b1;
      zz_rom_31[47] = 1'b1;
      zz_rom_31[48] = 1'b1;
      zz_rom_31[49] = 1'b1;
      zz_rom_31[50] = 1'b1;
      zz_rom_31[51] = 1'b1;
      zz_rom_31[52] = 1'b1;
      zz_rom_31[53] = 1'b1;
      zz_rom_31[54] = 1'b1;
      zz_rom_31[55] = 1'b1;
      zz_rom_31[56] = 1'b1;
      zz_rom_31[57] = 1'b1;
      zz_rom_31[58] = 1'b1;
      zz_rom_31[59] = 1'b1;
      zz_rom_31[60] = 1'b1;
      zz_rom_31[61] = 1'b1;
      zz_rom_31[62] = 1'b1;
      zz_rom_31[63] = 1'b1;
      zz_rom_31[64] = 1'b1;
      zz_rom_31[65] = 1'b1;
      zz_rom_31[66] = 1'b1;
      zz_rom_31[67] = 1'b1;
      zz_rom_31[68] = 1'b1;
      zz_rom_31[69] = 1'b1;
      zz_rom_31[70] = 1'b1;
      zz_rom_31[71] = 1'b1;
      zz_rom_31[72] = 1'b1;
      zz_rom_31[73] = 1'b1;
      zz_rom_31[74] = 1'b1;
      zz_rom_31[75] = 1'b1;
      zz_rom_31[76] = 1'b1;
      zz_rom_31[77] = 1'b1;
      zz_rom_31[78] = 1'b1;
      zz_rom_31[79] = 1'b1;
      zz_rom_31[80] = 1'b1;
      zz_rom_31[81] = 1'b1;
      zz_rom_31[82] = 1'b1;
      zz_rom_31[83] = 1'b1;
      zz_rom_31[84] = 1'b1;
      zz_rom_31[85] = 1'b1;
      zz_rom_31[86] = 1'b1;
      zz_rom_31[87] = 1'b1;
      zz_rom_31[88] = 1'b1;
      zz_rom_31[89] = 1'b1;
      zz_rom_31[90] = 1'b1;
      zz_rom_31[91] = 1'b1;
      zz_rom_31[92] = 1'b1;
      zz_rom_31[93] = 1'b1;
      zz_rom_31[94] = 1'b1;
      zz_rom_31[95] = 1'b1;
      zz_rom_31[96] = 1'b1;
      zz_rom_31[97] = 1'b0;
      zz_rom_31[98] = 1'b0;
      zz_rom_31[99] = 1'b0;
    end
  endfunction
  wire [99:0] _zz_32;
  function [99:0] zz_rom_32(input dummy);
    begin
      zz_rom_32[0] = 1'b0;
      zz_rom_32[1] = 1'b0;
      zz_rom_32[2] = 1'b0;
      zz_rom_32[3] = 1'b0;
      zz_rom_32[4] = 1'b1;
      zz_rom_32[5] = 1'b1;
      zz_rom_32[6] = 1'b1;
      zz_rom_32[7] = 1'b1;
      zz_rom_32[8] = 1'b1;
      zz_rom_32[9] = 1'b1;
      zz_rom_32[10] = 1'b1;
      zz_rom_32[11] = 1'b1;
      zz_rom_32[12] = 1'b1;
      zz_rom_32[13] = 1'b1;
      zz_rom_32[14] = 1'b1;
      zz_rom_32[15] = 1'b1;
      zz_rom_32[16] = 1'b1;
      zz_rom_32[17] = 1'b1;
      zz_rom_32[18] = 1'b1;
      zz_rom_32[19] = 1'b1;
      zz_rom_32[20] = 1'b1;
      zz_rom_32[21] = 1'b1;
      zz_rom_32[22] = 1'b1;
      zz_rom_32[23] = 1'b1;
      zz_rom_32[24] = 1'b1;
      zz_rom_32[25] = 1'b1;
      zz_rom_32[26] = 1'b1;
      zz_rom_32[27] = 1'b1;
      zz_rom_32[28] = 1'b1;
      zz_rom_32[29] = 1'b1;
      zz_rom_32[30] = 1'b1;
      zz_rom_32[31] = 1'b1;
      zz_rom_32[32] = 1'b1;
      zz_rom_32[33] = 1'b1;
      zz_rom_32[34] = 1'b1;
      zz_rom_32[35] = 1'b1;
      zz_rom_32[36] = 1'b1;
      zz_rom_32[37] = 1'b1;
      zz_rom_32[38] = 1'b1;
      zz_rom_32[39] = 1'b1;
      zz_rom_32[40] = 1'b1;
      zz_rom_32[41] = 1'b1;
      zz_rom_32[42] = 1'b1;
      zz_rom_32[43] = 1'b1;
      zz_rom_32[44] = 1'b1;
      zz_rom_32[45] = 1'b1;
      zz_rom_32[46] = 1'b1;
      zz_rom_32[47] = 1'b1;
      zz_rom_32[48] = 1'b1;
      zz_rom_32[49] = 1'b1;
      zz_rom_32[50] = 1'b1;
      zz_rom_32[51] = 1'b1;
      zz_rom_32[52] = 1'b1;
      zz_rom_32[53] = 1'b1;
      zz_rom_32[54] = 1'b1;
      zz_rom_32[55] = 1'b1;
      zz_rom_32[56] = 1'b1;
      zz_rom_32[57] = 1'b1;
      zz_rom_32[58] = 1'b1;
      zz_rom_32[59] = 1'b1;
      zz_rom_32[60] = 1'b1;
      zz_rom_32[61] = 1'b1;
      zz_rom_32[62] = 1'b1;
      zz_rom_32[63] = 1'b1;
      zz_rom_32[64] = 1'b1;
      zz_rom_32[65] = 1'b1;
      zz_rom_32[66] = 1'b1;
      zz_rom_32[67] = 1'b1;
      zz_rom_32[68] = 1'b1;
      zz_rom_32[69] = 1'b1;
      zz_rom_32[70] = 1'b1;
      zz_rom_32[71] = 1'b1;
      zz_rom_32[72] = 1'b1;
      zz_rom_32[73] = 1'b1;
      zz_rom_32[74] = 1'b1;
      zz_rom_32[75] = 1'b1;
      zz_rom_32[76] = 1'b1;
      zz_rom_32[77] = 1'b1;
      zz_rom_32[78] = 1'b1;
      zz_rom_32[79] = 1'b1;
      zz_rom_32[80] = 1'b1;
      zz_rom_32[81] = 1'b1;
      zz_rom_32[82] = 1'b1;
      zz_rom_32[83] = 1'b1;
      zz_rom_32[84] = 1'b1;
      zz_rom_32[85] = 1'b1;
      zz_rom_32[86] = 1'b1;
      zz_rom_32[87] = 1'b1;
      zz_rom_32[88] = 1'b1;
      zz_rom_32[89] = 1'b1;
      zz_rom_32[90] = 1'b1;
      zz_rom_32[91] = 1'b1;
      zz_rom_32[92] = 1'b1;
      zz_rom_32[93] = 1'b1;
      zz_rom_32[94] = 1'b1;
      zz_rom_32[95] = 1'b1;
      zz_rom_32[96] = 1'b1;
      zz_rom_32[97] = 1'b0;
      zz_rom_32[98] = 1'b0;
      zz_rom_32[99] = 1'b0;
    end
  endfunction
  wire [99:0] _zz_33;
  function [99:0] zz_rom_33(input dummy);
    begin
      zz_rom_33[0] = 1'b0;
      zz_rom_33[1] = 1'b0;
      zz_rom_33[2] = 1'b0;
      zz_rom_33[3] = 1'b1;
      zz_rom_33[4] = 1'b1;
      zz_rom_33[5] = 1'b1;
      zz_rom_33[6] = 1'b1;
      zz_rom_33[7] = 1'b1;
      zz_rom_33[8] = 1'b1;
      zz_rom_33[9] = 1'b1;
      zz_rom_33[10] = 1'b1;
      zz_rom_33[11] = 1'b1;
      zz_rom_33[12] = 1'b1;
      zz_rom_33[13] = 1'b1;
      zz_rom_33[14] = 1'b1;
      zz_rom_33[15] = 1'b1;
      zz_rom_33[16] = 1'b1;
      zz_rom_33[17] = 1'b1;
      zz_rom_33[18] = 1'b1;
      zz_rom_33[19] = 1'b1;
      zz_rom_33[20] = 1'b1;
      zz_rom_33[21] = 1'b1;
      zz_rom_33[22] = 1'b1;
      zz_rom_33[23] = 1'b1;
      zz_rom_33[24] = 1'b1;
      zz_rom_33[25] = 1'b1;
      zz_rom_33[26] = 1'b1;
      zz_rom_33[27] = 1'b1;
      zz_rom_33[28] = 1'b1;
      zz_rom_33[29] = 1'b1;
      zz_rom_33[30] = 1'b1;
      zz_rom_33[31] = 1'b1;
      zz_rom_33[32] = 1'b1;
      zz_rom_33[33] = 1'b1;
      zz_rom_33[34] = 1'b1;
      zz_rom_33[35] = 1'b1;
      zz_rom_33[36] = 1'b1;
      zz_rom_33[37] = 1'b1;
      zz_rom_33[38] = 1'b1;
      zz_rom_33[39] = 1'b1;
      zz_rom_33[40] = 1'b1;
      zz_rom_33[41] = 1'b1;
      zz_rom_33[42] = 1'b1;
      zz_rom_33[43] = 1'b1;
      zz_rom_33[44] = 1'b1;
      zz_rom_33[45] = 1'b1;
      zz_rom_33[46] = 1'b1;
      zz_rom_33[47] = 1'b1;
      zz_rom_33[48] = 1'b1;
      zz_rom_33[49] = 1'b1;
      zz_rom_33[50] = 1'b1;
      zz_rom_33[51] = 1'b1;
      zz_rom_33[52] = 1'b1;
      zz_rom_33[53] = 1'b1;
      zz_rom_33[54] = 1'b1;
      zz_rom_33[55] = 1'b1;
      zz_rom_33[56] = 1'b1;
      zz_rom_33[57] = 1'b1;
      zz_rom_33[58] = 1'b1;
      zz_rom_33[59] = 1'b1;
      zz_rom_33[60] = 1'b1;
      zz_rom_33[61] = 1'b1;
      zz_rom_33[62] = 1'b1;
      zz_rom_33[63] = 1'b1;
      zz_rom_33[64] = 1'b1;
      zz_rom_33[65] = 1'b1;
      zz_rom_33[66] = 1'b1;
      zz_rom_33[67] = 1'b1;
      zz_rom_33[68] = 1'b1;
      zz_rom_33[69] = 1'b1;
      zz_rom_33[70] = 1'b1;
      zz_rom_33[71] = 1'b1;
      zz_rom_33[72] = 1'b1;
      zz_rom_33[73] = 1'b1;
      zz_rom_33[74] = 1'b1;
      zz_rom_33[75] = 1'b1;
      zz_rom_33[76] = 1'b1;
      zz_rom_33[77] = 1'b1;
      zz_rom_33[78] = 1'b1;
      zz_rom_33[79] = 1'b1;
      zz_rom_33[80] = 1'b1;
      zz_rom_33[81] = 1'b1;
      zz_rom_33[82] = 1'b1;
      zz_rom_33[83] = 1'b1;
      zz_rom_33[84] = 1'b1;
      zz_rom_33[85] = 1'b1;
      zz_rom_33[86] = 1'b1;
      zz_rom_33[87] = 1'b1;
      zz_rom_33[88] = 1'b1;
      zz_rom_33[89] = 1'b1;
      zz_rom_33[90] = 1'b1;
      zz_rom_33[91] = 1'b1;
      zz_rom_33[92] = 1'b1;
      zz_rom_33[93] = 1'b1;
      zz_rom_33[94] = 1'b1;
      zz_rom_33[95] = 1'b1;
      zz_rom_33[96] = 1'b1;
      zz_rom_33[97] = 1'b1;
      zz_rom_33[98] = 1'b0;
      zz_rom_33[99] = 1'b0;
    end
  endfunction
  wire [99:0] _zz_34;
  function [99:0] zz_rom_34(input dummy);
    begin
      zz_rom_34[0] = 1'b0;
      zz_rom_34[1] = 1'b0;
      zz_rom_34[2] = 1'b0;
      zz_rom_34[3] = 1'b1;
      zz_rom_34[4] = 1'b1;
      zz_rom_34[5] = 1'b1;
      zz_rom_34[6] = 1'b1;
      zz_rom_34[7] = 1'b1;
      zz_rom_34[8] = 1'b1;
      zz_rom_34[9] = 1'b1;
      zz_rom_34[10] = 1'b1;
      zz_rom_34[11] = 1'b1;
      zz_rom_34[12] = 1'b1;
      zz_rom_34[13] = 1'b1;
      zz_rom_34[14] = 1'b1;
      zz_rom_34[15] = 1'b1;
      zz_rom_34[16] = 1'b1;
      zz_rom_34[17] = 1'b1;
      zz_rom_34[18] = 1'b1;
      zz_rom_34[19] = 1'b1;
      zz_rom_34[20] = 1'b1;
      zz_rom_34[21] = 1'b1;
      zz_rom_34[22] = 1'b1;
      zz_rom_34[23] = 1'b1;
      zz_rom_34[24] = 1'b1;
      zz_rom_34[25] = 1'b1;
      zz_rom_34[26] = 1'b1;
      zz_rom_34[27] = 1'b1;
      zz_rom_34[28] = 1'b1;
      zz_rom_34[29] = 1'b1;
      zz_rom_34[30] = 1'b1;
      zz_rom_34[31] = 1'b1;
      zz_rom_34[32] = 1'b1;
      zz_rom_34[33] = 1'b1;
      zz_rom_34[34] = 1'b1;
      zz_rom_34[35] = 1'b1;
      zz_rom_34[36] = 1'b1;
      zz_rom_34[37] = 1'b1;
      zz_rom_34[38] = 1'b1;
      zz_rom_34[39] = 1'b1;
      zz_rom_34[40] = 1'b1;
      zz_rom_34[41] = 1'b1;
      zz_rom_34[42] = 1'b1;
      zz_rom_34[43] = 1'b1;
      zz_rom_34[44] = 1'b1;
      zz_rom_34[45] = 1'b1;
      zz_rom_34[46] = 1'b1;
      zz_rom_34[47] = 1'b1;
      zz_rom_34[48] = 1'b1;
      zz_rom_34[49] = 1'b1;
      zz_rom_34[50] = 1'b1;
      zz_rom_34[51] = 1'b1;
      zz_rom_34[52] = 1'b1;
      zz_rom_34[53] = 1'b1;
      zz_rom_34[54] = 1'b1;
      zz_rom_34[55] = 1'b1;
      zz_rom_34[56] = 1'b1;
      zz_rom_34[57] = 1'b1;
      zz_rom_34[58] = 1'b1;
      zz_rom_34[59] = 1'b1;
      zz_rom_34[60] = 1'b1;
      zz_rom_34[61] = 1'b1;
      zz_rom_34[62] = 1'b1;
      zz_rom_34[63] = 1'b1;
      zz_rom_34[64] = 1'b1;
      zz_rom_34[65] = 1'b1;
      zz_rom_34[66] = 1'b1;
      zz_rom_34[67] = 1'b1;
      zz_rom_34[68] = 1'b1;
      zz_rom_34[69] = 1'b1;
      zz_rom_34[70] = 1'b1;
      zz_rom_34[71] = 1'b1;
      zz_rom_34[72] = 1'b1;
      zz_rom_34[73] = 1'b1;
      zz_rom_34[74] = 1'b1;
      zz_rom_34[75] = 1'b1;
      zz_rom_34[76] = 1'b1;
      zz_rom_34[77] = 1'b1;
      zz_rom_34[78] = 1'b1;
      zz_rom_34[79] = 1'b1;
      zz_rom_34[80] = 1'b1;
      zz_rom_34[81] = 1'b1;
      zz_rom_34[82] = 1'b1;
      zz_rom_34[83] = 1'b1;
      zz_rom_34[84] = 1'b1;
      zz_rom_34[85] = 1'b1;
      zz_rom_34[86] = 1'b1;
      zz_rom_34[87] = 1'b1;
      zz_rom_34[88] = 1'b1;
      zz_rom_34[89] = 1'b1;
      zz_rom_34[90] = 1'b1;
      zz_rom_34[91] = 1'b1;
      zz_rom_34[92] = 1'b1;
      zz_rom_34[93] = 1'b1;
      zz_rom_34[94] = 1'b1;
      zz_rom_34[95] = 1'b1;
      zz_rom_34[96] = 1'b1;
      zz_rom_34[97] = 1'b1;
      zz_rom_34[98] = 1'b0;
      zz_rom_34[99] = 1'b0;
    end
  endfunction
  wire [99:0] _zz_35;
  function [99:0] zz_rom_35(input dummy);
    begin
      zz_rom_35[0] = 1'b0;
      zz_rom_35[1] = 1'b0;
      zz_rom_35[2] = 1'b0;
      zz_rom_35[3] = 1'b1;
      zz_rom_35[4] = 1'b1;
      zz_rom_35[5] = 1'b1;
      zz_rom_35[6] = 1'b1;
      zz_rom_35[7] = 1'b1;
      zz_rom_35[8] = 1'b1;
      zz_rom_35[9] = 1'b1;
      zz_rom_35[10] = 1'b1;
      zz_rom_35[11] = 1'b1;
      zz_rom_35[12] = 1'b1;
      zz_rom_35[13] = 1'b1;
      zz_rom_35[14] = 1'b1;
      zz_rom_35[15] = 1'b1;
      zz_rom_35[16] = 1'b1;
      zz_rom_35[17] = 1'b1;
      zz_rom_35[18] = 1'b1;
      zz_rom_35[19] = 1'b1;
      zz_rom_35[20] = 1'b1;
      zz_rom_35[21] = 1'b1;
      zz_rom_35[22] = 1'b1;
      zz_rom_35[23] = 1'b1;
      zz_rom_35[24] = 1'b1;
      zz_rom_35[25] = 1'b1;
      zz_rom_35[26] = 1'b1;
      zz_rom_35[27] = 1'b1;
      zz_rom_35[28] = 1'b1;
      zz_rom_35[29] = 1'b1;
      zz_rom_35[30] = 1'b1;
      zz_rom_35[31] = 1'b1;
      zz_rom_35[32] = 1'b1;
      zz_rom_35[33] = 1'b1;
      zz_rom_35[34] = 1'b1;
      zz_rom_35[35] = 1'b1;
      zz_rom_35[36] = 1'b1;
      zz_rom_35[37] = 1'b1;
      zz_rom_35[38] = 1'b1;
      zz_rom_35[39] = 1'b1;
      zz_rom_35[40] = 1'b1;
      zz_rom_35[41] = 1'b1;
      zz_rom_35[42] = 1'b1;
      zz_rom_35[43] = 1'b1;
      zz_rom_35[44] = 1'b1;
      zz_rom_35[45] = 1'b1;
      zz_rom_35[46] = 1'b1;
      zz_rom_35[47] = 1'b1;
      zz_rom_35[48] = 1'b1;
      zz_rom_35[49] = 1'b1;
      zz_rom_35[50] = 1'b1;
      zz_rom_35[51] = 1'b1;
      zz_rom_35[52] = 1'b1;
      zz_rom_35[53] = 1'b1;
      zz_rom_35[54] = 1'b1;
      zz_rom_35[55] = 1'b1;
      zz_rom_35[56] = 1'b1;
      zz_rom_35[57] = 1'b1;
      zz_rom_35[58] = 1'b1;
      zz_rom_35[59] = 1'b1;
      zz_rom_35[60] = 1'b1;
      zz_rom_35[61] = 1'b1;
      zz_rom_35[62] = 1'b1;
      zz_rom_35[63] = 1'b1;
      zz_rom_35[64] = 1'b1;
      zz_rom_35[65] = 1'b1;
      zz_rom_35[66] = 1'b1;
      zz_rom_35[67] = 1'b1;
      zz_rom_35[68] = 1'b1;
      zz_rom_35[69] = 1'b1;
      zz_rom_35[70] = 1'b1;
      zz_rom_35[71] = 1'b1;
      zz_rom_35[72] = 1'b1;
      zz_rom_35[73] = 1'b1;
      zz_rom_35[74] = 1'b1;
      zz_rom_35[75] = 1'b1;
      zz_rom_35[76] = 1'b1;
      zz_rom_35[77] = 1'b1;
      zz_rom_35[78] = 1'b1;
      zz_rom_35[79] = 1'b1;
      zz_rom_35[80] = 1'b1;
      zz_rom_35[81] = 1'b1;
      zz_rom_35[82] = 1'b1;
      zz_rom_35[83] = 1'b1;
      zz_rom_35[84] = 1'b1;
      zz_rom_35[85] = 1'b1;
      zz_rom_35[86] = 1'b1;
      zz_rom_35[87] = 1'b1;
      zz_rom_35[88] = 1'b1;
      zz_rom_35[89] = 1'b1;
      zz_rom_35[90] = 1'b1;
      zz_rom_35[91] = 1'b1;
      zz_rom_35[92] = 1'b1;
      zz_rom_35[93] = 1'b1;
      zz_rom_35[94] = 1'b1;
      zz_rom_35[95] = 1'b1;
      zz_rom_35[96] = 1'b1;
      zz_rom_35[97] = 1'b1;
      zz_rom_35[98] = 1'b0;
      zz_rom_35[99] = 1'b0;
    end
  endfunction
  wire [99:0] _zz_36;
  function [99:0] zz_rom_36(input dummy);
    begin
      zz_rom_36[0] = 1'b0;
      zz_rom_36[1] = 1'b0;
      zz_rom_36[2] = 1'b1;
      zz_rom_36[3] = 1'b1;
      zz_rom_36[4] = 1'b1;
      zz_rom_36[5] = 1'b1;
      zz_rom_36[6] = 1'b1;
      zz_rom_36[7] = 1'b1;
      zz_rom_36[8] = 1'b1;
      zz_rom_36[9] = 1'b1;
      zz_rom_36[10] = 1'b1;
      zz_rom_36[11] = 1'b1;
      zz_rom_36[12] = 1'b1;
      zz_rom_36[13] = 1'b1;
      zz_rom_36[14] = 1'b1;
      zz_rom_36[15] = 1'b1;
      zz_rom_36[16] = 1'b1;
      zz_rom_36[17] = 1'b1;
      zz_rom_36[18] = 1'b1;
      zz_rom_36[19] = 1'b1;
      zz_rom_36[20] = 1'b1;
      zz_rom_36[21] = 1'b1;
      zz_rom_36[22] = 1'b1;
      zz_rom_36[23] = 1'b1;
      zz_rom_36[24] = 1'b1;
      zz_rom_36[25] = 1'b1;
      zz_rom_36[26] = 1'b1;
      zz_rom_36[27] = 1'b1;
      zz_rom_36[28] = 1'b1;
      zz_rom_36[29] = 1'b1;
      zz_rom_36[30] = 1'b1;
      zz_rom_36[31] = 1'b1;
      zz_rom_36[32] = 1'b1;
      zz_rom_36[33] = 1'b1;
      zz_rom_36[34] = 1'b1;
      zz_rom_36[35] = 1'b1;
      zz_rom_36[36] = 1'b1;
      zz_rom_36[37] = 1'b1;
      zz_rom_36[38] = 1'b1;
      zz_rom_36[39] = 1'b1;
      zz_rom_36[40] = 1'b1;
      zz_rom_36[41] = 1'b1;
      zz_rom_36[42] = 1'b1;
      zz_rom_36[43] = 1'b1;
      zz_rom_36[44] = 1'b1;
      zz_rom_36[45] = 1'b1;
      zz_rom_36[46] = 1'b1;
      zz_rom_36[47] = 1'b1;
      zz_rom_36[48] = 1'b1;
      zz_rom_36[49] = 1'b1;
      zz_rom_36[50] = 1'b1;
      zz_rom_36[51] = 1'b1;
      zz_rom_36[52] = 1'b1;
      zz_rom_36[53] = 1'b1;
      zz_rom_36[54] = 1'b1;
      zz_rom_36[55] = 1'b1;
      zz_rom_36[56] = 1'b1;
      zz_rom_36[57] = 1'b1;
      zz_rom_36[58] = 1'b1;
      zz_rom_36[59] = 1'b1;
      zz_rom_36[60] = 1'b1;
      zz_rom_36[61] = 1'b1;
      zz_rom_36[62] = 1'b1;
      zz_rom_36[63] = 1'b1;
      zz_rom_36[64] = 1'b1;
      zz_rom_36[65] = 1'b1;
      zz_rom_36[66] = 1'b1;
      zz_rom_36[67] = 1'b1;
      zz_rom_36[68] = 1'b1;
      zz_rom_36[69] = 1'b1;
      zz_rom_36[70] = 1'b1;
      zz_rom_36[71] = 1'b1;
      zz_rom_36[72] = 1'b1;
      zz_rom_36[73] = 1'b1;
      zz_rom_36[74] = 1'b1;
      zz_rom_36[75] = 1'b1;
      zz_rom_36[76] = 1'b1;
      zz_rom_36[77] = 1'b1;
      zz_rom_36[78] = 1'b1;
      zz_rom_36[79] = 1'b1;
      zz_rom_36[80] = 1'b1;
      zz_rom_36[81] = 1'b1;
      zz_rom_36[82] = 1'b1;
      zz_rom_36[83] = 1'b1;
      zz_rom_36[84] = 1'b1;
      zz_rom_36[85] = 1'b1;
      zz_rom_36[86] = 1'b1;
      zz_rom_36[87] = 1'b1;
      zz_rom_36[88] = 1'b1;
      zz_rom_36[89] = 1'b1;
      zz_rom_36[90] = 1'b1;
      zz_rom_36[91] = 1'b1;
      zz_rom_36[92] = 1'b1;
      zz_rom_36[93] = 1'b1;
      zz_rom_36[94] = 1'b1;
      zz_rom_36[95] = 1'b1;
      zz_rom_36[96] = 1'b1;
      zz_rom_36[97] = 1'b1;
      zz_rom_36[98] = 1'b1;
      zz_rom_36[99] = 1'b0;
    end
  endfunction
  wire [99:0] _zz_37;
  function [99:0] zz_rom_37(input dummy);
    begin
      zz_rom_37[0] = 1'b0;
      zz_rom_37[1] = 1'b0;
      zz_rom_37[2] = 1'b1;
      zz_rom_37[3] = 1'b1;
      zz_rom_37[4] = 1'b1;
      zz_rom_37[5] = 1'b1;
      zz_rom_37[6] = 1'b1;
      zz_rom_37[7] = 1'b1;
      zz_rom_37[8] = 1'b1;
      zz_rom_37[9] = 1'b1;
      zz_rom_37[10] = 1'b1;
      zz_rom_37[11] = 1'b1;
      zz_rom_37[12] = 1'b1;
      zz_rom_37[13] = 1'b1;
      zz_rom_37[14] = 1'b1;
      zz_rom_37[15] = 1'b1;
      zz_rom_37[16] = 1'b1;
      zz_rom_37[17] = 1'b1;
      zz_rom_37[18] = 1'b1;
      zz_rom_37[19] = 1'b1;
      zz_rom_37[20] = 1'b1;
      zz_rom_37[21] = 1'b1;
      zz_rom_37[22] = 1'b1;
      zz_rom_37[23] = 1'b1;
      zz_rom_37[24] = 1'b1;
      zz_rom_37[25] = 1'b1;
      zz_rom_37[26] = 1'b1;
      zz_rom_37[27] = 1'b1;
      zz_rom_37[28] = 1'b1;
      zz_rom_37[29] = 1'b1;
      zz_rom_37[30] = 1'b1;
      zz_rom_37[31] = 1'b1;
      zz_rom_37[32] = 1'b1;
      zz_rom_37[33] = 1'b1;
      zz_rom_37[34] = 1'b1;
      zz_rom_37[35] = 1'b1;
      zz_rom_37[36] = 1'b1;
      zz_rom_37[37] = 1'b1;
      zz_rom_37[38] = 1'b1;
      zz_rom_37[39] = 1'b1;
      zz_rom_37[40] = 1'b1;
      zz_rom_37[41] = 1'b1;
      zz_rom_37[42] = 1'b1;
      zz_rom_37[43] = 1'b1;
      zz_rom_37[44] = 1'b1;
      zz_rom_37[45] = 1'b1;
      zz_rom_37[46] = 1'b1;
      zz_rom_37[47] = 1'b1;
      zz_rom_37[48] = 1'b1;
      zz_rom_37[49] = 1'b1;
      zz_rom_37[50] = 1'b1;
      zz_rom_37[51] = 1'b1;
      zz_rom_37[52] = 1'b1;
      zz_rom_37[53] = 1'b1;
      zz_rom_37[54] = 1'b1;
      zz_rom_37[55] = 1'b1;
      zz_rom_37[56] = 1'b1;
      zz_rom_37[57] = 1'b1;
      zz_rom_37[58] = 1'b1;
      zz_rom_37[59] = 1'b1;
      zz_rom_37[60] = 1'b1;
      zz_rom_37[61] = 1'b1;
      zz_rom_37[62] = 1'b1;
      zz_rom_37[63] = 1'b1;
      zz_rom_37[64] = 1'b1;
      zz_rom_37[65] = 1'b1;
      zz_rom_37[66] = 1'b1;
      zz_rom_37[67] = 1'b1;
      zz_rom_37[68] = 1'b1;
      zz_rom_37[69] = 1'b1;
      zz_rom_37[70] = 1'b1;
      zz_rom_37[71] = 1'b1;
      zz_rom_37[72] = 1'b1;
      zz_rom_37[73] = 1'b1;
      zz_rom_37[74] = 1'b1;
      zz_rom_37[75] = 1'b1;
      zz_rom_37[76] = 1'b1;
      zz_rom_37[77] = 1'b1;
      zz_rom_37[78] = 1'b1;
      zz_rom_37[79] = 1'b1;
      zz_rom_37[80] = 1'b1;
      zz_rom_37[81] = 1'b1;
      zz_rom_37[82] = 1'b1;
      zz_rom_37[83] = 1'b1;
      zz_rom_37[84] = 1'b1;
      zz_rom_37[85] = 1'b1;
      zz_rom_37[86] = 1'b1;
      zz_rom_37[87] = 1'b1;
      zz_rom_37[88] = 1'b1;
      zz_rom_37[89] = 1'b1;
      zz_rom_37[90] = 1'b1;
      zz_rom_37[91] = 1'b1;
      zz_rom_37[92] = 1'b1;
      zz_rom_37[93] = 1'b1;
      zz_rom_37[94] = 1'b1;
      zz_rom_37[95] = 1'b1;
      zz_rom_37[96] = 1'b1;
      zz_rom_37[97] = 1'b1;
      zz_rom_37[98] = 1'b1;
      zz_rom_37[99] = 1'b0;
    end
  endfunction
  wire [99:0] _zz_38;
  function [99:0] zz_rom_38(input dummy);
    begin
      zz_rom_38[0] = 1'b0;
      zz_rom_38[1] = 1'b0;
      zz_rom_38[2] = 1'b1;
      zz_rom_38[3] = 1'b1;
      zz_rom_38[4] = 1'b1;
      zz_rom_38[5] = 1'b1;
      zz_rom_38[6] = 1'b1;
      zz_rom_38[7] = 1'b1;
      zz_rom_38[8] = 1'b1;
      zz_rom_38[9] = 1'b1;
      zz_rom_38[10] = 1'b1;
      zz_rom_38[11] = 1'b1;
      zz_rom_38[12] = 1'b1;
      zz_rom_38[13] = 1'b1;
      zz_rom_38[14] = 1'b1;
      zz_rom_38[15] = 1'b1;
      zz_rom_38[16] = 1'b1;
      zz_rom_38[17] = 1'b1;
      zz_rom_38[18] = 1'b1;
      zz_rom_38[19] = 1'b1;
      zz_rom_38[20] = 1'b1;
      zz_rom_38[21] = 1'b1;
      zz_rom_38[22] = 1'b1;
      zz_rom_38[23] = 1'b1;
      zz_rom_38[24] = 1'b1;
      zz_rom_38[25] = 1'b1;
      zz_rom_38[26] = 1'b1;
      zz_rom_38[27] = 1'b1;
      zz_rom_38[28] = 1'b1;
      zz_rom_38[29] = 1'b1;
      zz_rom_38[30] = 1'b1;
      zz_rom_38[31] = 1'b1;
      zz_rom_38[32] = 1'b1;
      zz_rom_38[33] = 1'b1;
      zz_rom_38[34] = 1'b1;
      zz_rom_38[35] = 1'b1;
      zz_rom_38[36] = 1'b1;
      zz_rom_38[37] = 1'b1;
      zz_rom_38[38] = 1'b1;
      zz_rom_38[39] = 1'b1;
      zz_rom_38[40] = 1'b1;
      zz_rom_38[41] = 1'b1;
      zz_rom_38[42] = 1'b1;
      zz_rom_38[43] = 1'b1;
      zz_rom_38[44] = 1'b1;
      zz_rom_38[45] = 1'b1;
      zz_rom_38[46] = 1'b1;
      zz_rom_38[47] = 1'b1;
      zz_rom_38[48] = 1'b1;
      zz_rom_38[49] = 1'b1;
      zz_rom_38[50] = 1'b1;
      zz_rom_38[51] = 1'b1;
      zz_rom_38[52] = 1'b1;
      zz_rom_38[53] = 1'b1;
      zz_rom_38[54] = 1'b1;
      zz_rom_38[55] = 1'b1;
      zz_rom_38[56] = 1'b1;
      zz_rom_38[57] = 1'b1;
      zz_rom_38[58] = 1'b1;
      zz_rom_38[59] = 1'b1;
      zz_rom_38[60] = 1'b1;
      zz_rom_38[61] = 1'b1;
      zz_rom_38[62] = 1'b1;
      zz_rom_38[63] = 1'b1;
      zz_rom_38[64] = 1'b1;
      zz_rom_38[65] = 1'b1;
      zz_rom_38[66] = 1'b1;
      zz_rom_38[67] = 1'b1;
      zz_rom_38[68] = 1'b1;
      zz_rom_38[69] = 1'b1;
      zz_rom_38[70] = 1'b1;
      zz_rom_38[71] = 1'b1;
      zz_rom_38[72] = 1'b1;
      zz_rom_38[73] = 1'b1;
      zz_rom_38[74] = 1'b1;
      zz_rom_38[75] = 1'b1;
      zz_rom_38[76] = 1'b1;
      zz_rom_38[77] = 1'b1;
      zz_rom_38[78] = 1'b1;
      zz_rom_38[79] = 1'b1;
      zz_rom_38[80] = 1'b1;
      zz_rom_38[81] = 1'b1;
      zz_rom_38[82] = 1'b1;
      zz_rom_38[83] = 1'b1;
      zz_rom_38[84] = 1'b1;
      zz_rom_38[85] = 1'b1;
      zz_rom_38[86] = 1'b1;
      zz_rom_38[87] = 1'b1;
      zz_rom_38[88] = 1'b1;
      zz_rom_38[89] = 1'b1;
      zz_rom_38[90] = 1'b1;
      zz_rom_38[91] = 1'b1;
      zz_rom_38[92] = 1'b1;
      zz_rom_38[93] = 1'b1;
      zz_rom_38[94] = 1'b1;
      zz_rom_38[95] = 1'b1;
      zz_rom_38[96] = 1'b1;
      zz_rom_38[97] = 1'b1;
      zz_rom_38[98] = 1'b1;
      zz_rom_38[99] = 1'b0;
    end
  endfunction
  wire [99:0] _zz_39;
  function [99:0] zz_rom_39(input dummy);
    begin
      zz_rom_39[0] = 1'b0;
      zz_rom_39[1] = 1'b0;
      zz_rom_39[2] = 1'b1;
      zz_rom_39[3] = 1'b1;
      zz_rom_39[4] = 1'b1;
      zz_rom_39[5] = 1'b1;
      zz_rom_39[6] = 1'b1;
      zz_rom_39[7] = 1'b1;
      zz_rom_39[8] = 1'b1;
      zz_rom_39[9] = 1'b1;
      zz_rom_39[10] = 1'b1;
      zz_rom_39[11] = 1'b1;
      zz_rom_39[12] = 1'b1;
      zz_rom_39[13] = 1'b1;
      zz_rom_39[14] = 1'b1;
      zz_rom_39[15] = 1'b1;
      zz_rom_39[16] = 1'b1;
      zz_rom_39[17] = 1'b1;
      zz_rom_39[18] = 1'b1;
      zz_rom_39[19] = 1'b1;
      zz_rom_39[20] = 1'b1;
      zz_rom_39[21] = 1'b1;
      zz_rom_39[22] = 1'b1;
      zz_rom_39[23] = 1'b1;
      zz_rom_39[24] = 1'b1;
      zz_rom_39[25] = 1'b1;
      zz_rom_39[26] = 1'b1;
      zz_rom_39[27] = 1'b1;
      zz_rom_39[28] = 1'b1;
      zz_rom_39[29] = 1'b1;
      zz_rom_39[30] = 1'b1;
      zz_rom_39[31] = 1'b1;
      zz_rom_39[32] = 1'b1;
      zz_rom_39[33] = 1'b1;
      zz_rom_39[34] = 1'b1;
      zz_rom_39[35] = 1'b1;
      zz_rom_39[36] = 1'b1;
      zz_rom_39[37] = 1'b1;
      zz_rom_39[38] = 1'b1;
      zz_rom_39[39] = 1'b1;
      zz_rom_39[40] = 1'b1;
      zz_rom_39[41] = 1'b1;
      zz_rom_39[42] = 1'b1;
      zz_rom_39[43] = 1'b1;
      zz_rom_39[44] = 1'b1;
      zz_rom_39[45] = 1'b1;
      zz_rom_39[46] = 1'b1;
      zz_rom_39[47] = 1'b1;
      zz_rom_39[48] = 1'b1;
      zz_rom_39[49] = 1'b1;
      zz_rom_39[50] = 1'b1;
      zz_rom_39[51] = 1'b1;
      zz_rom_39[52] = 1'b1;
      zz_rom_39[53] = 1'b1;
      zz_rom_39[54] = 1'b1;
      zz_rom_39[55] = 1'b1;
      zz_rom_39[56] = 1'b1;
      zz_rom_39[57] = 1'b1;
      zz_rom_39[58] = 1'b1;
      zz_rom_39[59] = 1'b1;
      zz_rom_39[60] = 1'b1;
      zz_rom_39[61] = 1'b1;
      zz_rom_39[62] = 1'b1;
      zz_rom_39[63] = 1'b1;
      zz_rom_39[64] = 1'b1;
      zz_rom_39[65] = 1'b1;
      zz_rom_39[66] = 1'b1;
      zz_rom_39[67] = 1'b1;
      zz_rom_39[68] = 1'b1;
      zz_rom_39[69] = 1'b1;
      zz_rom_39[70] = 1'b1;
      zz_rom_39[71] = 1'b1;
      zz_rom_39[72] = 1'b1;
      zz_rom_39[73] = 1'b1;
      zz_rom_39[74] = 1'b1;
      zz_rom_39[75] = 1'b1;
      zz_rom_39[76] = 1'b1;
      zz_rom_39[77] = 1'b1;
      zz_rom_39[78] = 1'b1;
      zz_rom_39[79] = 1'b1;
      zz_rom_39[80] = 1'b1;
      zz_rom_39[81] = 1'b1;
      zz_rom_39[82] = 1'b1;
      zz_rom_39[83] = 1'b1;
      zz_rom_39[84] = 1'b1;
      zz_rom_39[85] = 1'b1;
      zz_rom_39[86] = 1'b1;
      zz_rom_39[87] = 1'b1;
      zz_rom_39[88] = 1'b1;
      zz_rom_39[89] = 1'b1;
      zz_rom_39[90] = 1'b1;
      zz_rom_39[91] = 1'b1;
      zz_rom_39[92] = 1'b1;
      zz_rom_39[93] = 1'b1;
      zz_rom_39[94] = 1'b1;
      zz_rom_39[95] = 1'b1;
      zz_rom_39[96] = 1'b1;
      zz_rom_39[97] = 1'b1;
      zz_rom_39[98] = 1'b1;
      zz_rom_39[99] = 1'b0;
    end
  endfunction
  wire [99:0] _zz_40;
  function [99:0] zz_rom_40(input dummy);
    begin
      zz_rom_40[0] = 1'b0;
      zz_rom_40[1] = 1'b0;
      zz_rom_40[2] = 1'b1;
      zz_rom_40[3] = 1'b1;
      zz_rom_40[4] = 1'b1;
      zz_rom_40[5] = 1'b1;
      zz_rom_40[6] = 1'b1;
      zz_rom_40[7] = 1'b1;
      zz_rom_40[8] = 1'b1;
      zz_rom_40[9] = 1'b1;
      zz_rom_40[10] = 1'b1;
      zz_rom_40[11] = 1'b1;
      zz_rom_40[12] = 1'b1;
      zz_rom_40[13] = 1'b1;
      zz_rom_40[14] = 1'b1;
      zz_rom_40[15] = 1'b1;
      zz_rom_40[16] = 1'b1;
      zz_rom_40[17] = 1'b1;
      zz_rom_40[18] = 1'b1;
      zz_rom_40[19] = 1'b1;
      zz_rom_40[20] = 1'b1;
      zz_rom_40[21] = 1'b1;
      zz_rom_40[22] = 1'b1;
      zz_rom_40[23] = 1'b1;
      zz_rom_40[24] = 1'b1;
      zz_rom_40[25] = 1'b1;
      zz_rom_40[26] = 1'b1;
      zz_rom_40[27] = 1'b1;
      zz_rom_40[28] = 1'b1;
      zz_rom_40[29] = 1'b1;
      zz_rom_40[30] = 1'b1;
      zz_rom_40[31] = 1'b1;
      zz_rom_40[32] = 1'b1;
      zz_rom_40[33] = 1'b1;
      zz_rom_40[34] = 1'b1;
      zz_rom_40[35] = 1'b1;
      zz_rom_40[36] = 1'b1;
      zz_rom_40[37] = 1'b1;
      zz_rom_40[38] = 1'b1;
      zz_rom_40[39] = 1'b1;
      zz_rom_40[40] = 1'b1;
      zz_rom_40[41] = 1'b1;
      zz_rom_40[42] = 1'b1;
      zz_rom_40[43] = 1'b1;
      zz_rom_40[44] = 1'b1;
      zz_rom_40[45] = 1'b1;
      zz_rom_40[46] = 1'b1;
      zz_rom_40[47] = 1'b1;
      zz_rom_40[48] = 1'b1;
      zz_rom_40[49] = 1'b1;
      zz_rom_40[50] = 1'b1;
      zz_rom_40[51] = 1'b1;
      zz_rom_40[52] = 1'b1;
      zz_rom_40[53] = 1'b1;
      zz_rom_40[54] = 1'b1;
      zz_rom_40[55] = 1'b1;
      zz_rom_40[56] = 1'b1;
      zz_rom_40[57] = 1'b1;
      zz_rom_40[58] = 1'b1;
      zz_rom_40[59] = 1'b1;
      zz_rom_40[60] = 1'b1;
      zz_rom_40[61] = 1'b1;
      zz_rom_40[62] = 1'b1;
      zz_rom_40[63] = 1'b1;
      zz_rom_40[64] = 1'b1;
      zz_rom_40[65] = 1'b1;
      zz_rom_40[66] = 1'b1;
      zz_rom_40[67] = 1'b1;
      zz_rom_40[68] = 1'b1;
      zz_rom_40[69] = 1'b1;
      zz_rom_40[70] = 1'b1;
      zz_rom_40[71] = 1'b1;
      zz_rom_40[72] = 1'b1;
      zz_rom_40[73] = 1'b1;
      zz_rom_40[74] = 1'b1;
      zz_rom_40[75] = 1'b1;
      zz_rom_40[76] = 1'b1;
      zz_rom_40[77] = 1'b1;
      zz_rom_40[78] = 1'b1;
      zz_rom_40[79] = 1'b1;
      zz_rom_40[80] = 1'b1;
      zz_rom_40[81] = 1'b1;
      zz_rom_40[82] = 1'b1;
      zz_rom_40[83] = 1'b1;
      zz_rom_40[84] = 1'b1;
      zz_rom_40[85] = 1'b1;
      zz_rom_40[86] = 1'b1;
      zz_rom_40[87] = 1'b1;
      zz_rom_40[88] = 1'b1;
      zz_rom_40[89] = 1'b1;
      zz_rom_40[90] = 1'b1;
      zz_rom_40[91] = 1'b1;
      zz_rom_40[92] = 1'b1;
      zz_rom_40[93] = 1'b1;
      zz_rom_40[94] = 1'b1;
      zz_rom_40[95] = 1'b1;
      zz_rom_40[96] = 1'b1;
      zz_rom_40[97] = 1'b1;
      zz_rom_40[98] = 1'b1;
      zz_rom_40[99] = 1'b0;
    end
  endfunction
  wire [99:0] _zz_41;
  function [99:0] zz_rom_41(input dummy);
    begin
      zz_rom_41[0] = 1'b0;
      zz_rom_41[1] = 1'b1;
      zz_rom_41[2] = 1'b1;
      zz_rom_41[3] = 1'b1;
      zz_rom_41[4] = 1'b1;
      zz_rom_41[5] = 1'b1;
      zz_rom_41[6] = 1'b1;
      zz_rom_41[7] = 1'b1;
      zz_rom_41[8] = 1'b1;
      zz_rom_41[9] = 1'b1;
      zz_rom_41[10] = 1'b1;
      zz_rom_41[11] = 1'b1;
      zz_rom_41[12] = 1'b1;
      zz_rom_41[13] = 1'b1;
      zz_rom_41[14] = 1'b1;
      zz_rom_41[15] = 1'b1;
      zz_rom_41[16] = 1'b1;
      zz_rom_41[17] = 1'b1;
      zz_rom_41[18] = 1'b1;
      zz_rom_41[19] = 1'b1;
      zz_rom_41[20] = 1'b1;
      zz_rom_41[21] = 1'b1;
      zz_rom_41[22] = 1'b1;
      zz_rom_41[23] = 1'b1;
      zz_rom_41[24] = 1'b1;
      zz_rom_41[25] = 1'b1;
      zz_rom_41[26] = 1'b1;
      zz_rom_41[27] = 1'b1;
      zz_rom_41[28] = 1'b1;
      zz_rom_41[29] = 1'b1;
      zz_rom_41[30] = 1'b1;
      zz_rom_41[31] = 1'b1;
      zz_rom_41[32] = 1'b1;
      zz_rom_41[33] = 1'b1;
      zz_rom_41[34] = 1'b1;
      zz_rom_41[35] = 1'b1;
      zz_rom_41[36] = 1'b1;
      zz_rom_41[37] = 1'b1;
      zz_rom_41[38] = 1'b1;
      zz_rom_41[39] = 1'b1;
      zz_rom_41[40] = 1'b1;
      zz_rom_41[41] = 1'b1;
      zz_rom_41[42] = 1'b1;
      zz_rom_41[43] = 1'b1;
      zz_rom_41[44] = 1'b1;
      zz_rom_41[45] = 1'b1;
      zz_rom_41[46] = 1'b1;
      zz_rom_41[47] = 1'b1;
      zz_rom_41[48] = 1'b1;
      zz_rom_41[49] = 1'b1;
      zz_rom_41[50] = 1'b1;
      zz_rom_41[51] = 1'b1;
      zz_rom_41[52] = 1'b1;
      zz_rom_41[53] = 1'b1;
      zz_rom_41[54] = 1'b1;
      zz_rom_41[55] = 1'b1;
      zz_rom_41[56] = 1'b1;
      zz_rom_41[57] = 1'b1;
      zz_rom_41[58] = 1'b1;
      zz_rom_41[59] = 1'b1;
      zz_rom_41[60] = 1'b1;
      zz_rom_41[61] = 1'b1;
      zz_rom_41[62] = 1'b1;
      zz_rom_41[63] = 1'b1;
      zz_rom_41[64] = 1'b1;
      zz_rom_41[65] = 1'b1;
      zz_rom_41[66] = 1'b1;
      zz_rom_41[67] = 1'b1;
      zz_rom_41[68] = 1'b1;
      zz_rom_41[69] = 1'b1;
      zz_rom_41[70] = 1'b1;
      zz_rom_41[71] = 1'b1;
      zz_rom_41[72] = 1'b1;
      zz_rom_41[73] = 1'b1;
      zz_rom_41[74] = 1'b1;
      zz_rom_41[75] = 1'b1;
      zz_rom_41[76] = 1'b1;
      zz_rom_41[77] = 1'b1;
      zz_rom_41[78] = 1'b1;
      zz_rom_41[79] = 1'b1;
      zz_rom_41[80] = 1'b1;
      zz_rom_41[81] = 1'b1;
      zz_rom_41[82] = 1'b1;
      zz_rom_41[83] = 1'b1;
      zz_rom_41[84] = 1'b1;
      zz_rom_41[85] = 1'b1;
      zz_rom_41[86] = 1'b1;
      zz_rom_41[87] = 1'b1;
      zz_rom_41[88] = 1'b1;
      zz_rom_41[89] = 1'b1;
      zz_rom_41[90] = 1'b1;
      zz_rom_41[91] = 1'b1;
      zz_rom_41[92] = 1'b1;
      zz_rom_41[93] = 1'b1;
      zz_rom_41[94] = 1'b1;
      zz_rom_41[95] = 1'b1;
      zz_rom_41[96] = 1'b1;
      zz_rom_41[97] = 1'b1;
      zz_rom_41[98] = 1'b1;
      zz_rom_41[99] = 1'b1;
    end
  endfunction
  wire [99:0] _zz_42;
  function [99:0] zz_rom_42(input dummy);
    begin
      zz_rom_42[0] = 1'b0;
      zz_rom_42[1] = 1'b1;
      zz_rom_42[2] = 1'b1;
      zz_rom_42[3] = 1'b1;
      zz_rom_42[4] = 1'b1;
      zz_rom_42[5] = 1'b1;
      zz_rom_42[6] = 1'b1;
      zz_rom_42[7] = 1'b1;
      zz_rom_42[8] = 1'b1;
      zz_rom_42[9] = 1'b1;
      zz_rom_42[10] = 1'b1;
      zz_rom_42[11] = 1'b1;
      zz_rom_42[12] = 1'b1;
      zz_rom_42[13] = 1'b1;
      zz_rom_42[14] = 1'b1;
      zz_rom_42[15] = 1'b1;
      zz_rom_42[16] = 1'b1;
      zz_rom_42[17] = 1'b1;
      zz_rom_42[18] = 1'b1;
      zz_rom_42[19] = 1'b1;
      zz_rom_42[20] = 1'b1;
      zz_rom_42[21] = 1'b1;
      zz_rom_42[22] = 1'b1;
      zz_rom_42[23] = 1'b1;
      zz_rom_42[24] = 1'b1;
      zz_rom_42[25] = 1'b1;
      zz_rom_42[26] = 1'b1;
      zz_rom_42[27] = 1'b1;
      zz_rom_42[28] = 1'b1;
      zz_rom_42[29] = 1'b1;
      zz_rom_42[30] = 1'b1;
      zz_rom_42[31] = 1'b1;
      zz_rom_42[32] = 1'b1;
      zz_rom_42[33] = 1'b1;
      zz_rom_42[34] = 1'b1;
      zz_rom_42[35] = 1'b1;
      zz_rom_42[36] = 1'b1;
      zz_rom_42[37] = 1'b1;
      zz_rom_42[38] = 1'b1;
      zz_rom_42[39] = 1'b1;
      zz_rom_42[40] = 1'b1;
      zz_rom_42[41] = 1'b1;
      zz_rom_42[42] = 1'b1;
      zz_rom_42[43] = 1'b1;
      zz_rom_42[44] = 1'b1;
      zz_rom_42[45] = 1'b1;
      zz_rom_42[46] = 1'b1;
      zz_rom_42[47] = 1'b1;
      zz_rom_42[48] = 1'b1;
      zz_rom_42[49] = 1'b1;
      zz_rom_42[50] = 1'b1;
      zz_rom_42[51] = 1'b1;
      zz_rom_42[52] = 1'b1;
      zz_rom_42[53] = 1'b1;
      zz_rom_42[54] = 1'b1;
      zz_rom_42[55] = 1'b1;
      zz_rom_42[56] = 1'b1;
      zz_rom_42[57] = 1'b1;
      zz_rom_42[58] = 1'b1;
      zz_rom_42[59] = 1'b1;
      zz_rom_42[60] = 1'b1;
      zz_rom_42[61] = 1'b1;
      zz_rom_42[62] = 1'b1;
      zz_rom_42[63] = 1'b1;
      zz_rom_42[64] = 1'b1;
      zz_rom_42[65] = 1'b1;
      zz_rom_42[66] = 1'b1;
      zz_rom_42[67] = 1'b1;
      zz_rom_42[68] = 1'b1;
      zz_rom_42[69] = 1'b1;
      zz_rom_42[70] = 1'b1;
      zz_rom_42[71] = 1'b1;
      zz_rom_42[72] = 1'b1;
      zz_rom_42[73] = 1'b1;
      zz_rom_42[74] = 1'b1;
      zz_rom_42[75] = 1'b1;
      zz_rom_42[76] = 1'b1;
      zz_rom_42[77] = 1'b1;
      zz_rom_42[78] = 1'b1;
      zz_rom_42[79] = 1'b1;
      zz_rom_42[80] = 1'b1;
      zz_rom_42[81] = 1'b1;
      zz_rom_42[82] = 1'b1;
      zz_rom_42[83] = 1'b1;
      zz_rom_42[84] = 1'b1;
      zz_rom_42[85] = 1'b1;
      zz_rom_42[86] = 1'b1;
      zz_rom_42[87] = 1'b1;
      zz_rom_42[88] = 1'b1;
      zz_rom_42[89] = 1'b1;
      zz_rom_42[90] = 1'b1;
      zz_rom_42[91] = 1'b1;
      zz_rom_42[92] = 1'b1;
      zz_rom_42[93] = 1'b1;
      zz_rom_42[94] = 1'b1;
      zz_rom_42[95] = 1'b1;
      zz_rom_42[96] = 1'b1;
      zz_rom_42[97] = 1'b1;
      zz_rom_42[98] = 1'b1;
      zz_rom_42[99] = 1'b1;
    end
  endfunction
  wire [99:0] _zz_43;
  function [99:0] zz_rom_43(input dummy);
    begin
      zz_rom_43[0] = 1'b0;
      zz_rom_43[1] = 1'b1;
      zz_rom_43[2] = 1'b1;
      zz_rom_43[3] = 1'b1;
      zz_rom_43[4] = 1'b1;
      zz_rom_43[5] = 1'b1;
      zz_rom_43[6] = 1'b1;
      zz_rom_43[7] = 1'b1;
      zz_rom_43[8] = 1'b1;
      zz_rom_43[9] = 1'b1;
      zz_rom_43[10] = 1'b1;
      zz_rom_43[11] = 1'b1;
      zz_rom_43[12] = 1'b1;
      zz_rom_43[13] = 1'b1;
      zz_rom_43[14] = 1'b1;
      zz_rom_43[15] = 1'b1;
      zz_rom_43[16] = 1'b1;
      zz_rom_43[17] = 1'b1;
      zz_rom_43[18] = 1'b1;
      zz_rom_43[19] = 1'b1;
      zz_rom_43[20] = 1'b1;
      zz_rom_43[21] = 1'b1;
      zz_rom_43[22] = 1'b1;
      zz_rom_43[23] = 1'b1;
      zz_rom_43[24] = 1'b1;
      zz_rom_43[25] = 1'b1;
      zz_rom_43[26] = 1'b1;
      zz_rom_43[27] = 1'b1;
      zz_rom_43[28] = 1'b1;
      zz_rom_43[29] = 1'b1;
      zz_rom_43[30] = 1'b1;
      zz_rom_43[31] = 1'b1;
      zz_rom_43[32] = 1'b1;
      zz_rom_43[33] = 1'b1;
      zz_rom_43[34] = 1'b1;
      zz_rom_43[35] = 1'b1;
      zz_rom_43[36] = 1'b1;
      zz_rom_43[37] = 1'b1;
      zz_rom_43[38] = 1'b1;
      zz_rom_43[39] = 1'b1;
      zz_rom_43[40] = 1'b1;
      zz_rom_43[41] = 1'b1;
      zz_rom_43[42] = 1'b1;
      zz_rom_43[43] = 1'b1;
      zz_rom_43[44] = 1'b1;
      zz_rom_43[45] = 1'b1;
      zz_rom_43[46] = 1'b1;
      zz_rom_43[47] = 1'b1;
      zz_rom_43[48] = 1'b1;
      zz_rom_43[49] = 1'b1;
      zz_rom_43[50] = 1'b1;
      zz_rom_43[51] = 1'b1;
      zz_rom_43[52] = 1'b1;
      zz_rom_43[53] = 1'b1;
      zz_rom_43[54] = 1'b1;
      zz_rom_43[55] = 1'b1;
      zz_rom_43[56] = 1'b1;
      zz_rom_43[57] = 1'b1;
      zz_rom_43[58] = 1'b1;
      zz_rom_43[59] = 1'b1;
      zz_rom_43[60] = 1'b1;
      zz_rom_43[61] = 1'b1;
      zz_rom_43[62] = 1'b1;
      zz_rom_43[63] = 1'b1;
      zz_rom_43[64] = 1'b1;
      zz_rom_43[65] = 1'b1;
      zz_rom_43[66] = 1'b1;
      zz_rom_43[67] = 1'b1;
      zz_rom_43[68] = 1'b1;
      zz_rom_43[69] = 1'b1;
      zz_rom_43[70] = 1'b1;
      zz_rom_43[71] = 1'b1;
      zz_rom_43[72] = 1'b1;
      zz_rom_43[73] = 1'b1;
      zz_rom_43[74] = 1'b1;
      zz_rom_43[75] = 1'b1;
      zz_rom_43[76] = 1'b1;
      zz_rom_43[77] = 1'b1;
      zz_rom_43[78] = 1'b1;
      zz_rom_43[79] = 1'b1;
      zz_rom_43[80] = 1'b1;
      zz_rom_43[81] = 1'b1;
      zz_rom_43[82] = 1'b1;
      zz_rom_43[83] = 1'b1;
      zz_rom_43[84] = 1'b1;
      zz_rom_43[85] = 1'b1;
      zz_rom_43[86] = 1'b1;
      zz_rom_43[87] = 1'b1;
      zz_rom_43[88] = 1'b1;
      zz_rom_43[89] = 1'b1;
      zz_rom_43[90] = 1'b1;
      zz_rom_43[91] = 1'b1;
      zz_rom_43[92] = 1'b1;
      zz_rom_43[93] = 1'b1;
      zz_rom_43[94] = 1'b1;
      zz_rom_43[95] = 1'b1;
      zz_rom_43[96] = 1'b1;
      zz_rom_43[97] = 1'b1;
      zz_rom_43[98] = 1'b1;
      zz_rom_43[99] = 1'b1;
    end
  endfunction
  wire [99:0] _zz_44;
  function [99:0] zz_rom_44(input dummy);
    begin
      zz_rom_44[0] = 1'b0;
      zz_rom_44[1] = 1'b1;
      zz_rom_44[2] = 1'b1;
      zz_rom_44[3] = 1'b1;
      zz_rom_44[4] = 1'b1;
      zz_rom_44[5] = 1'b1;
      zz_rom_44[6] = 1'b1;
      zz_rom_44[7] = 1'b1;
      zz_rom_44[8] = 1'b1;
      zz_rom_44[9] = 1'b1;
      zz_rom_44[10] = 1'b1;
      zz_rom_44[11] = 1'b1;
      zz_rom_44[12] = 1'b1;
      zz_rom_44[13] = 1'b1;
      zz_rom_44[14] = 1'b1;
      zz_rom_44[15] = 1'b1;
      zz_rom_44[16] = 1'b1;
      zz_rom_44[17] = 1'b1;
      zz_rom_44[18] = 1'b1;
      zz_rom_44[19] = 1'b1;
      zz_rom_44[20] = 1'b1;
      zz_rom_44[21] = 1'b1;
      zz_rom_44[22] = 1'b1;
      zz_rom_44[23] = 1'b1;
      zz_rom_44[24] = 1'b1;
      zz_rom_44[25] = 1'b1;
      zz_rom_44[26] = 1'b1;
      zz_rom_44[27] = 1'b1;
      zz_rom_44[28] = 1'b1;
      zz_rom_44[29] = 1'b1;
      zz_rom_44[30] = 1'b1;
      zz_rom_44[31] = 1'b1;
      zz_rom_44[32] = 1'b1;
      zz_rom_44[33] = 1'b1;
      zz_rom_44[34] = 1'b1;
      zz_rom_44[35] = 1'b1;
      zz_rom_44[36] = 1'b1;
      zz_rom_44[37] = 1'b1;
      zz_rom_44[38] = 1'b1;
      zz_rom_44[39] = 1'b1;
      zz_rom_44[40] = 1'b1;
      zz_rom_44[41] = 1'b1;
      zz_rom_44[42] = 1'b1;
      zz_rom_44[43] = 1'b1;
      zz_rom_44[44] = 1'b1;
      zz_rom_44[45] = 1'b1;
      zz_rom_44[46] = 1'b1;
      zz_rom_44[47] = 1'b1;
      zz_rom_44[48] = 1'b1;
      zz_rom_44[49] = 1'b1;
      zz_rom_44[50] = 1'b1;
      zz_rom_44[51] = 1'b1;
      zz_rom_44[52] = 1'b1;
      zz_rom_44[53] = 1'b1;
      zz_rom_44[54] = 1'b1;
      zz_rom_44[55] = 1'b1;
      zz_rom_44[56] = 1'b1;
      zz_rom_44[57] = 1'b1;
      zz_rom_44[58] = 1'b1;
      zz_rom_44[59] = 1'b1;
      zz_rom_44[60] = 1'b1;
      zz_rom_44[61] = 1'b1;
      zz_rom_44[62] = 1'b1;
      zz_rom_44[63] = 1'b1;
      zz_rom_44[64] = 1'b1;
      zz_rom_44[65] = 1'b1;
      zz_rom_44[66] = 1'b1;
      zz_rom_44[67] = 1'b1;
      zz_rom_44[68] = 1'b1;
      zz_rom_44[69] = 1'b1;
      zz_rom_44[70] = 1'b1;
      zz_rom_44[71] = 1'b1;
      zz_rom_44[72] = 1'b1;
      zz_rom_44[73] = 1'b1;
      zz_rom_44[74] = 1'b1;
      zz_rom_44[75] = 1'b1;
      zz_rom_44[76] = 1'b1;
      zz_rom_44[77] = 1'b1;
      zz_rom_44[78] = 1'b1;
      zz_rom_44[79] = 1'b1;
      zz_rom_44[80] = 1'b1;
      zz_rom_44[81] = 1'b1;
      zz_rom_44[82] = 1'b1;
      zz_rom_44[83] = 1'b1;
      zz_rom_44[84] = 1'b1;
      zz_rom_44[85] = 1'b1;
      zz_rom_44[86] = 1'b1;
      zz_rom_44[87] = 1'b1;
      zz_rom_44[88] = 1'b1;
      zz_rom_44[89] = 1'b1;
      zz_rom_44[90] = 1'b1;
      zz_rom_44[91] = 1'b1;
      zz_rom_44[92] = 1'b1;
      zz_rom_44[93] = 1'b1;
      zz_rom_44[94] = 1'b1;
      zz_rom_44[95] = 1'b1;
      zz_rom_44[96] = 1'b1;
      zz_rom_44[97] = 1'b1;
      zz_rom_44[98] = 1'b1;
      zz_rom_44[99] = 1'b1;
    end
  endfunction
  wire [99:0] _zz_45;
  function [99:0] zz_rom_45(input dummy);
    begin
      zz_rom_45[0] = 1'b0;
      zz_rom_45[1] = 1'b1;
      zz_rom_45[2] = 1'b1;
      zz_rom_45[3] = 1'b1;
      zz_rom_45[4] = 1'b1;
      zz_rom_45[5] = 1'b1;
      zz_rom_45[6] = 1'b1;
      zz_rom_45[7] = 1'b1;
      zz_rom_45[8] = 1'b1;
      zz_rom_45[9] = 1'b1;
      zz_rom_45[10] = 1'b1;
      zz_rom_45[11] = 1'b1;
      zz_rom_45[12] = 1'b1;
      zz_rom_45[13] = 1'b1;
      zz_rom_45[14] = 1'b1;
      zz_rom_45[15] = 1'b1;
      zz_rom_45[16] = 1'b1;
      zz_rom_45[17] = 1'b1;
      zz_rom_45[18] = 1'b1;
      zz_rom_45[19] = 1'b1;
      zz_rom_45[20] = 1'b1;
      zz_rom_45[21] = 1'b1;
      zz_rom_45[22] = 1'b1;
      zz_rom_45[23] = 1'b1;
      zz_rom_45[24] = 1'b1;
      zz_rom_45[25] = 1'b1;
      zz_rom_45[26] = 1'b1;
      zz_rom_45[27] = 1'b1;
      zz_rom_45[28] = 1'b1;
      zz_rom_45[29] = 1'b1;
      zz_rom_45[30] = 1'b1;
      zz_rom_45[31] = 1'b1;
      zz_rom_45[32] = 1'b1;
      zz_rom_45[33] = 1'b1;
      zz_rom_45[34] = 1'b1;
      zz_rom_45[35] = 1'b1;
      zz_rom_45[36] = 1'b1;
      zz_rom_45[37] = 1'b1;
      zz_rom_45[38] = 1'b1;
      zz_rom_45[39] = 1'b1;
      zz_rom_45[40] = 1'b1;
      zz_rom_45[41] = 1'b1;
      zz_rom_45[42] = 1'b1;
      zz_rom_45[43] = 1'b1;
      zz_rom_45[44] = 1'b1;
      zz_rom_45[45] = 1'b1;
      zz_rom_45[46] = 1'b1;
      zz_rom_45[47] = 1'b1;
      zz_rom_45[48] = 1'b1;
      zz_rom_45[49] = 1'b1;
      zz_rom_45[50] = 1'b1;
      zz_rom_45[51] = 1'b1;
      zz_rom_45[52] = 1'b1;
      zz_rom_45[53] = 1'b1;
      zz_rom_45[54] = 1'b1;
      zz_rom_45[55] = 1'b1;
      zz_rom_45[56] = 1'b1;
      zz_rom_45[57] = 1'b1;
      zz_rom_45[58] = 1'b1;
      zz_rom_45[59] = 1'b1;
      zz_rom_45[60] = 1'b1;
      zz_rom_45[61] = 1'b1;
      zz_rom_45[62] = 1'b1;
      zz_rom_45[63] = 1'b1;
      zz_rom_45[64] = 1'b1;
      zz_rom_45[65] = 1'b1;
      zz_rom_45[66] = 1'b1;
      zz_rom_45[67] = 1'b1;
      zz_rom_45[68] = 1'b1;
      zz_rom_45[69] = 1'b1;
      zz_rom_45[70] = 1'b1;
      zz_rom_45[71] = 1'b1;
      zz_rom_45[72] = 1'b1;
      zz_rom_45[73] = 1'b1;
      zz_rom_45[74] = 1'b1;
      zz_rom_45[75] = 1'b1;
      zz_rom_45[76] = 1'b1;
      zz_rom_45[77] = 1'b1;
      zz_rom_45[78] = 1'b1;
      zz_rom_45[79] = 1'b1;
      zz_rom_45[80] = 1'b1;
      zz_rom_45[81] = 1'b1;
      zz_rom_45[82] = 1'b1;
      zz_rom_45[83] = 1'b1;
      zz_rom_45[84] = 1'b1;
      zz_rom_45[85] = 1'b1;
      zz_rom_45[86] = 1'b1;
      zz_rom_45[87] = 1'b1;
      zz_rom_45[88] = 1'b1;
      zz_rom_45[89] = 1'b1;
      zz_rom_45[90] = 1'b1;
      zz_rom_45[91] = 1'b1;
      zz_rom_45[92] = 1'b1;
      zz_rom_45[93] = 1'b1;
      zz_rom_45[94] = 1'b1;
      zz_rom_45[95] = 1'b1;
      zz_rom_45[96] = 1'b1;
      zz_rom_45[97] = 1'b1;
      zz_rom_45[98] = 1'b1;
      zz_rom_45[99] = 1'b1;
    end
  endfunction
  wire [99:0] _zz_46;
  function [99:0] zz_rom_46(input dummy);
    begin
      zz_rom_46[0] = 1'b0;
      zz_rom_46[1] = 1'b1;
      zz_rom_46[2] = 1'b1;
      zz_rom_46[3] = 1'b1;
      zz_rom_46[4] = 1'b1;
      zz_rom_46[5] = 1'b1;
      zz_rom_46[6] = 1'b1;
      zz_rom_46[7] = 1'b1;
      zz_rom_46[8] = 1'b1;
      zz_rom_46[9] = 1'b1;
      zz_rom_46[10] = 1'b1;
      zz_rom_46[11] = 1'b1;
      zz_rom_46[12] = 1'b1;
      zz_rom_46[13] = 1'b1;
      zz_rom_46[14] = 1'b1;
      zz_rom_46[15] = 1'b1;
      zz_rom_46[16] = 1'b1;
      zz_rom_46[17] = 1'b1;
      zz_rom_46[18] = 1'b1;
      zz_rom_46[19] = 1'b1;
      zz_rom_46[20] = 1'b1;
      zz_rom_46[21] = 1'b1;
      zz_rom_46[22] = 1'b1;
      zz_rom_46[23] = 1'b1;
      zz_rom_46[24] = 1'b1;
      zz_rom_46[25] = 1'b1;
      zz_rom_46[26] = 1'b1;
      zz_rom_46[27] = 1'b1;
      zz_rom_46[28] = 1'b1;
      zz_rom_46[29] = 1'b1;
      zz_rom_46[30] = 1'b1;
      zz_rom_46[31] = 1'b1;
      zz_rom_46[32] = 1'b1;
      zz_rom_46[33] = 1'b1;
      zz_rom_46[34] = 1'b1;
      zz_rom_46[35] = 1'b1;
      zz_rom_46[36] = 1'b1;
      zz_rom_46[37] = 1'b1;
      zz_rom_46[38] = 1'b1;
      zz_rom_46[39] = 1'b1;
      zz_rom_46[40] = 1'b1;
      zz_rom_46[41] = 1'b1;
      zz_rom_46[42] = 1'b1;
      zz_rom_46[43] = 1'b1;
      zz_rom_46[44] = 1'b1;
      zz_rom_46[45] = 1'b1;
      zz_rom_46[46] = 1'b1;
      zz_rom_46[47] = 1'b1;
      zz_rom_46[48] = 1'b1;
      zz_rom_46[49] = 1'b1;
      zz_rom_46[50] = 1'b1;
      zz_rom_46[51] = 1'b1;
      zz_rom_46[52] = 1'b1;
      zz_rom_46[53] = 1'b1;
      zz_rom_46[54] = 1'b1;
      zz_rom_46[55] = 1'b1;
      zz_rom_46[56] = 1'b1;
      zz_rom_46[57] = 1'b1;
      zz_rom_46[58] = 1'b1;
      zz_rom_46[59] = 1'b1;
      zz_rom_46[60] = 1'b1;
      zz_rom_46[61] = 1'b1;
      zz_rom_46[62] = 1'b1;
      zz_rom_46[63] = 1'b1;
      zz_rom_46[64] = 1'b1;
      zz_rom_46[65] = 1'b1;
      zz_rom_46[66] = 1'b1;
      zz_rom_46[67] = 1'b1;
      zz_rom_46[68] = 1'b1;
      zz_rom_46[69] = 1'b1;
      zz_rom_46[70] = 1'b1;
      zz_rom_46[71] = 1'b1;
      zz_rom_46[72] = 1'b1;
      zz_rom_46[73] = 1'b1;
      zz_rom_46[74] = 1'b1;
      zz_rom_46[75] = 1'b1;
      zz_rom_46[76] = 1'b1;
      zz_rom_46[77] = 1'b1;
      zz_rom_46[78] = 1'b1;
      zz_rom_46[79] = 1'b1;
      zz_rom_46[80] = 1'b1;
      zz_rom_46[81] = 1'b1;
      zz_rom_46[82] = 1'b1;
      zz_rom_46[83] = 1'b1;
      zz_rom_46[84] = 1'b1;
      zz_rom_46[85] = 1'b1;
      zz_rom_46[86] = 1'b1;
      zz_rom_46[87] = 1'b1;
      zz_rom_46[88] = 1'b1;
      zz_rom_46[89] = 1'b1;
      zz_rom_46[90] = 1'b1;
      zz_rom_46[91] = 1'b1;
      zz_rom_46[92] = 1'b1;
      zz_rom_46[93] = 1'b1;
      zz_rom_46[94] = 1'b1;
      zz_rom_46[95] = 1'b1;
      zz_rom_46[96] = 1'b1;
      zz_rom_46[97] = 1'b1;
      zz_rom_46[98] = 1'b1;
      zz_rom_46[99] = 1'b1;
    end
  endfunction
  wire [99:0] _zz_47;
  function [99:0] zz_rom_47(input dummy);
    begin
      zz_rom_47[0] = 1'b0;
      zz_rom_47[1] = 1'b1;
      zz_rom_47[2] = 1'b1;
      zz_rom_47[3] = 1'b1;
      zz_rom_47[4] = 1'b1;
      zz_rom_47[5] = 1'b1;
      zz_rom_47[6] = 1'b1;
      zz_rom_47[7] = 1'b1;
      zz_rom_47[8] = 1'b1;
      zz_rom_47[9] = 1'b1;
      zz_rom_47[10] = 1'b1;
      zz_rom_47[11] = 1'b1;
      zz_rom_47[12] = 1'b1;
      zz_rom_47[13] = 1'b1;
      zz_rom_47[14] = 1'b1;
      zz_rom_47[15] = 1'b1;
      zz_rom_47[16] = 1'b1;
      zz_rom_47[17] = 1'b1;
      zz_rom_47[18] = 1'b1;
      zz_rom_47[19] = 1'b1;
      zz_rom_47[20] = 1'b1;
      zz_rom_47[21] = 1'b1;
      zz_rom_47[22] = 1'b1;
      zz_rom_47[23] = 1'b1;
      zz_rom_47[24] = 1'b1;
      zz_rom_47[25] = 1'b1;
      zz_rom_47[26] = 1'b1;
      zz_rom_47[27] = 1'b1;
      zz_rom_47[28] = 1'b1;
      zz_rom_47[29] = 1'b1;
      zz_rom_47[30] = 1'b1;
      zz_rom_47[31] = 1'b1;
      zz_rom_47[32] = 1'b1;
      zz_rom_47[33] = 1'b1;
      zz_rom_47[34] = 1'b1;
      zz_rom_47[35] = 1'b1;
      zz_rom_47[36] = 1'b1;
      zz_rom_47[37] = 1'b1;
      zz_rom_47[38] = 1'b1;
      zz_rom_47[39] = 1'b1;
      zz_rom_47[40] = 1'b1;
      zz_rom_47[41] = 1'b1;
      zz_rom_47[42] = 1'b1;
      zz_rom_47[43] = 1'b1;
      zz_rom_47[44] = 1'b1;
      zz_rom_47[45] = 1'b1;
      zz_rom_47[46] = 1'b1;
      zz_rom_47[47] = 1'b1;
      zz_rom_47[48] = 1'b1;
      zz_rom_47[49] = 1'b1;
      zz_rom_47[50] = 1'b1;
      zz_rom_47[51] = 1'b1;
      zz_rom_47[52] = 1'b1;
      zz_rom_47[53] = 1'b1;
      zz_rom_47[54] = 1'b1;
      zz_rom_47[55] = 1'b1;
      zz_rom_47[56] = 1'b1;
      zz_rom_47[57] = 1'b1;
      zz_rom_47[58] = 1'b1;
      zz_rom_47[59] = 1'b1;
      zz_rom_47[60] = 1'b1;
      zz_rom_47[61] = 1'b1;
      zz_rom_47[62] = 1'b1;
      zz_rom_47[63] = 1'b1;
      zz_rom_47[64] = 1'b1;
      zz_rom_47[65] = 1'b1;
      zz_rom_47[66] = 1'b1;
      zz_rom_47[67] = 1'b1;
      zz_rom_47[68] = 1'b1;
      zz_rom_47[69] = 1'b1;
      zz_rom_47[70] = 1'b1;
      zz_rom_47[71] = 1'b1;
      zz_rom_47[72] = 1'b1;
      zz_rom_47[73] = 1'b1;
      zz_rom_47[74] = 1'b1;
      zz_rom_47[75] = 1'b1;
      zz_rom_47[76] = 1'b1;
      zz_rom_47[77] = 1'b1;
      zz_rom_47[78] = 1'b1;
      zz_rom_47[79] = 1'b1;
      zz_rom_47[80] = 1'b1;
      zz_rom_47[81] = 1'b1;
      zz_rom_47[82] = 1'b1;
      zz_rom_47[83] = 1'b1;
      zz_rom_47[84] = 1'b1;
      zz_rom_47[85] = 1'b1;
      zz_rom_47[86] = 1'b1;
      zz_rom_47[87] = 1'b1;
      zz_rom_47[88] = 1'b1;
      zz_rom_47[89] = 1'b1;
      zz_rom_47[90] = 1'b1;
      zz_rom_47[91] = 1'b1;
      zz_rom_47[92] = 1'b1;
      zz_rom_47[93] = 1'b1;
      zz_rom_47[94] = 1'b1;
      zz_rom_47[95] = 1'b1;
      zz_rom_47[96] = 1'b1;
      zz_rom_47[97] = 1'b1;
      zz_rom_47[98] = 1'b1;
      zz_rom_47[99] = 1'b1;
    end
  endfunction
  wire [99:0] _zz_48;
  function [99:0] zz_rom_48(input dummy);
    begin
      zz_rom_48[0] = 1'b0;
      zz_rom_48[1] = 1'b1;
      zz_rom_48[2] = 1'b1;
      zz_rom_48[3] = 1'b1;
      zz_rom_48[4] = 1'b1;
      zz_rom_48[5] = 1'b1;
      zz_rom_48[6] = 1'b1;
      zz_rom_48[7] = 1'b1;
      zz_rom_48[8] = 1'b1;
      zz_rom_48[9] = 1'b1;
      zz_rom_48[10] = 1'b1;
      zz_rom_48[11] = 1'b1;
      zz_rom_48[12] = 1'b1;
      zz_rom_48[13] = 1'b1;
      zz_rom_48[14] = 1'b1;
      zz_rom_48[15] = 1'b1;
      zz_rom_48[16] = 1'b1;
      zz_rom_48[17] = 1'b1;
      zz_rom_48[18] = 1'b1;
      zz_rom_48[19] = 1'b1;
      zz_rom_48[20] = 1'b1;
      zz_rom_48[21] = 1'b1;
      zz_rom_48[22] = 1'b1;
      zz_rom_48[23] = 1'b1;
      zz_rom_48[24] = 1'b1;
      zz_rom_48[25] = 1'b1;
      zz_rom_48[26] = 1'b1;
      zz_rom_48[27] = 1'b1;
      zz_rom_48[28] = 1'b1;
      zz_rom_48[29] = 1'b1;
      zz_rom_48[30] = 1'b1;
      zz_rom_48[31] = 1'b1;
      zz_rom_48[32] = 1'b1;
      zz_rom_48[33] = 1'b1;
      zz_rom_48[34] = 1'b1;
      zz_rom_48[35] = 1'b1;
      zz_rom_48[36] = 1'b1;
      zz_rom_48[37] = 1'b1;
      zz_rom_48[38] = 1'b1;
      zz_rom_48[39] = 1'b1;
      zz_rom_48[40] = 1'b1;
      zz_rom_48[41] = 1'b1;
      zz_rom_48[42] = 1'b1;
      zz_rom_48[43] = 1'b1;
      zz_rom_48[44] = 1'b1;
      zz_rom_48[45] = 1'b1;
      zz_rom_48[46] = 1'b1;
      zz_rom_48[47] = 1'b1;
      zz_rom_48[48] = 1'b1;
      zz_rom_48[49] = 1'b1;
      zz_rom_48[50] = 1'b1;
      zz_rom_48[51] = 1'b1;
      zz_rom_48[52] = 1'b1;
      zz_rom_48[53] = 1'b1;
      zz_rom_48[54] = 1'b1;
      zz_rom_48[55] = 1'b1;
      zz_rom_48[56] = 1'b1;
      zz_rom_48[57] = 1'b1;
      zz_rom_48[58] = 1'b1;
      zz_rom_48[59] = 1'b1;
      zz_rom_48[60] = 1'b1;
      zz_rom_48[61] = 1'b1;
      zz_rom_48[62] = 1'b1;
      zz_rom_48[63] = 1'b1;
      zz_rom_48[64] = 1'b1;
      zz_rom_48[65] = 1'b1;
      zz_rom_48[66] = 1'b1;
      zz_rom_48[67] = 1'b1;
      zz_rom_48[68] = 1'b1;
      zz_rom_48[69] = 1'b1;
      zz_rom_48[70] = 1'b1;
      zz_rom_48[71] = 1'b1;
      zz_rom_48[72] = 1'b1;
      zz_rom_48[73] = 1'b1;
      zz_rom_48[74] = 1'b1;
      zz_rom_48[75] = 1'b1;
      zz_rom_48[76] = 1'b1;
      zz_rom_48[77] = 1'b1;
      zz_rom_48[78] = 1'b1;
      zz_rom_48[79] = 1'b1;
      zz_rom_48[80] = 1'b1;
      zz_rom_48[81] = 1'b1;
      zz_rom_48[82] = 1'b1;
      zz_rom_48[83] = 1'b1;
      zz_rom_48[84] = 1'b1;
      zz_rom_48[85] = 1'b1;
      zz_rom_48[86] = 1'b1;
      zz_rom_48[87] = 1'b1;
      zz_rom_48[88] = 1'b1;
      zz_rom_48[89] = 1'b1;
      zz_rom_48[90] = 1'b1;
      zz_rom_48[91] = 1'b1;
      zz_rom_48[92] = 1'b1;
      zz_rom_48[93] = 1'b1;
      zz_rom_48[94] = 1'b1;
      zz_rom_48[95] = 1'b1;
      zz_rom_48[96] = 1'b1;
      zz_rom_48[97] = 1'b1;
      zz_rom_48[98] = 1'b1;
      zz_rom_48[99] = 1'b1;
    end
  endfunction
  wire [99:0] _zz_49;
  function [99:0] zz_rom_49(input dummy);
    begin
      zz_rom_49[0] = 1'b0;
      zz_rom_49[1] = 1'b1;
      zz_rom_49[2] = 1'b1;
      zz_rom_49[3] = 1'b1;
      zz_rom_49[4] = 1'b1;
      zz_rom_49[5] = 1'b1;
      zz_rom_49[6] = 1'b1;
      zz_rom_49[7] = 1'b1;
      zz_rom_49[8] = 1'b1;
      zz_rom_49[9] = 1'b1;
      zz_rom_49[10] = 1'b1;
      zz_rom_49[11] = 1'b1;
      zz_rom_49[12] = 1'b1;
      zz_rom_49[13] = 1'b1;
      zz_rom_49[14] = 1'b1;
      zz_rom_49[15] = 1'b1;
      zz_rom_49[16] = 1'b1;
      zz_rom_49[17] = 1'b1;
      zz_rom_49[18] = 1'b1;
      zz_rom_49[19] = 1'b1;
      zz_rom_49[20] = 1'b1;
      zz_rom_49[21] = 1'b1;
      zz_rom_49[22] = 1'b1;
      zz_rom_49[23] = 1'b1;
      zz_rom_49[24] = 1'b1;
      zz_rom_49[25] = 1'b1;
      zz_rom_49[26] = 1'b1;
      zz_rom_49[27] = 1'b1;
      zz_rom_49[28] = 1'b1;
      zz_rom_49[29] = 1'b1;
      zz_rom_49[30] = 1'b1;
      zz_rom_49[31] = 1'b1;
      zz_rom_49[32] = 1'b1;
      zz_rom_49[33] = 1'b1;
      zz_rom_49[34] = 1'b1;
      zz_rom_49[35] = 1'b1;
      zz_rom_49[36] = 1'b1;
      zz_rom_49[37] = 1'b1;
      zz_rom_49[38] = 1'b1;
      zz_rom_49[39] = 1'b1;
      zz_rom_49[40] = 1'b1;
      zz_rom_49[41] = 1'b1;
      zz_rom_49[42] = 1'b1;
      zz_rom_49[43] = 1'b1;
      zz_rom_49[44] = 1'b1;
      zz_rom_49[45] = 1'b1;
      zz_rom_49[46] = 1'b1;
      zz_rom_49[47] = 1'b1;
      zz_rom_49[48] = 1'b1;
      zz_rom_49[49] = 1'b1;
      zz_rom_49[50] = 1'b1;
      zz_rom_49[51] = 1'b1;
      zz_rom_49[52] = 1'b1;
      zz_rom_49[53] = 1'b1;
      zz_rom_49[54] = 1'b1;
      zz_rom_49[55] = 1'b1;
      zz_rom_49[56] = 1'b1;
      zz_rom_49[57] = 1'b1;
      zz_rom_49[58] = 1'b1;
      zz_rom_49[59] = 1'b1;
      zz_rom_49[60] = 1'b1;
      zz_rom_49[61] = 1'b1;
      zz_rom_49[62] = 1'b1;
      zz_rom_49[63] = 1'b1;
      zz_rom_49[64] = 1'b1;
      zz_rom_49[65] = 1'b1;
      zz_rom_49[66] = 1'b1;
      zz_rom_49[67] = 1'b1;
      zz_rom_49[68] = 1'b1;
      zz_rom_49[69] = 1'b1;
      zz_rom_49[70] = 1'b1;
      zz_rom_49[71] = 1'b1;
      zz_rom_49[72] = 1'b1;
      zz_rom_49[73] = 1'b1;
      zz_rom_49[74] = 1'b1;
      zz_rom_49[75] = 1'b1;
      zz_rom_49[76] = 1'b1;
      zz_rom_49[77] = 1'b1;
      zz_rom_49[78] = 1'b1;
      zz_rom_49[79] = 1'b1;
      zz_rom_49[80] = 1'b1;
      zz_rom_49[81] = 1'b1;
      zz_rom_49[82] = 1'b1;
      zz_rom_49[83] = 1'b1;
      zz_rom_49[84] = 1'b1;
      zz_rom_49[85] = 1'b1;
      zz_rom_49[86] = 1'b1;
      zz_rom_49[87] = 1'b1;
      zz_rom_49[88] = 1'b1;
      zz_rom_49[89] = 1'b1;
      zz_rom_49[90] = 1'b1;
      zz_rom_49[91] = 1'b1;
      zz_rom_49[92] = 1'b1;
      zz_rom_49[93] = 1'b1;
      zz_rom_49[94] = 1'b1;
      zz_rom_49[95] = 1'b1;
      zz_rom_49[96] = 1'b1;
      zz_rom_49[97] = 1'b1;
      zz_rom_49[98] = 1'b1;
      zz_rom_49[99] = 1'b1;
    end
  endfunction
  wire [99:0] _zz_50;
  function [99:0] zz_rom_50(input dummy);
    begin
      zz_rom_50[0] = 1'b1;
      zz_rom_50[1] = 1'b1;
      zz_rom_50[2] = 1'b1;
      zz_rom_50[3] = 1'b1;
      zz_rom_50[4] = 1'b1;
      zz_rom_50[5] = 1'b1;
      zz_rom_50[6] = 1'b1;
      zz_rom_50[7] = 1'b1;
      zz_rom_50[8] = 1'b1;
      zz_rom_50[9] = 1'b1;
      zz_rom_50[10] = 1'b1;
      zz_rom_50[11] = 1'b1;
      zz_rom_50[12] = 1'b1;
      zz_rom_50[13] = 1'b1;
      zz_rom_50[14] = 1'b1;
      zz_rom_50[15] = 1'b1;
      zz_rom_50[16] = 1'b1;
      zz_rom_50[17] = 1'b1;
      zz_rom_50[18] = 1'b1;
      zz_rom_50[19] = 1'b1;
      zz_rom_50[20] = 1'b1;
      zz_rom_50[21] = 1'b1;
      zz_rom_50[22] = 1'b1;
      zz_rom_50[23] = 1'b1;
      zz_rom_50[24] = 1'b1;
      zz_rom_50[25] = 1'b1;
      zz_rom_50[26] = 1'b1;
      zz_rom_50[27] = 1'b1;
      zz_rom_50[28] = 1'b1;
      zz_rom_50[29] = 1'b1;
      zz_rom_50[30] = 1'b1;
      zz_rom_50[31] = 1'b1;
      zz_rom_50[32] = 1'b1;
      zz_rom_50[33] = 1'b1;
      zz_rom_50[34] = 1'b1;
      zz_rom_50[35] = 1'b1;
      zz_rom_50[36] = 1'b1;
      zz_rom_50[37] = 1'b1;
      zz_rom_50[38] = 1'b1;
      zz_rom_50[39] = 1'b1;
      zz_rom_50[40] = 1'b1;
      zz_rom_50[41] = 1'b1;
      zz_rom_50[42] = 1'b1;
      zz_rom_50[43] = 1'b1;
      zz_rom_50[44] = 1'b1;
      zz_rom_50[45] = 1'b1;
      zz_rom_50[46] = 1'b1;
      zz_rom_50[47] = 1'b1;
      zz_rom_50[48] = 1'b1;
      zz_rom_50[49] = 1'b1;
      zz_rom_50[50] = 1'b1;
      zz_rom_50[51] = 1'b1;
      zz_rom_50[52] = 1'b1;
      zz_rom_50[53] = 1'b1;
      zz_rom_50[54] = 1'b1;
      zz_rom_50[55] = 1'b1;
      zz_rom_50[56] = 1'b1;
      zz_rom_50[57] = 1'b1;
      zz_rom_50[58] = 1'b1;
      zz_rom_50[59] = 1'b1;
      zz_rom_50[60] = 1'b1;
      zz_rom_50[61] = 1'b1;
      zz_rom_50[62] = 1'b1;
      zz_rom_50[63] = 1'b1;
      zz_rom_50[64] = 1'b1;
      zz_rom_50[65] = 1'b1;
      zz_rom_50[66] = 1'b1;
      zz_rom_50[67] = 1'b1;
      zz_rom_50[68] = 1'b1;
      zz_rom_50[69] = 1'b1;
      zz_rom_50[70] = 1'b1;
      zz_rom_50[71] = 1'b1;
      zz_rom_50[72] = 1'b1;
      zz_rom_50[73] = 1'b1;
      zz_rom_50[74] = 1'b1;
      zz_rom_50[75] = 1'b1;
      zz_rom_50[76] = 1'b1;
      zz_rom_50[77] = 1'b1;
      zz_rom_50[78] = 1'b1;
      zz_rom_50[79] = 1'b1;
      zz_rom_50[80] = 1'b1;
      zz_rom_50[81] = 1'b1;
      zz_rom_50[82] = 1'b1;
      zz_rom_50[83] = 1'b1;
      zz_rom_50[84] = 1'b1;
      zz_rom_50[85] = 1'b1;
      zz_rom_50[86] = 1'b1;
      zz_rom_50[87] = 1'b1;
      zz_rom_50[88] = 1'b1;
      zz_rom_50[89] = 1'b1;
      zz_rom_50[90] = 1'b1;
      zz_rom_50[91] = 1'b1;
      zz_rom_50[92] = 1'b1;
      zz_rom_50[93] = 1'b1;
      zz_rom_50[94] = 1'b1;
      zz_rom_50[95] = 1'b1;
      zz_rom_50[96] = 1'b1;
      zz_rom_50[97] = 1'b1;
      zz_rom_50[98] = 1'b1;
      zz_rom_50[99] = 1'b1;
    end
  endfunction
  wire [99:0] _zz_51;
  function [99:0] zz_rom_51(input dummy);
    begin
      zz_rom_51[0] = 1'b0;
      zz_rom_51[1] = 1'b1;
      zz_rom_51[2] = 1'b1;
      zz_rom_51[3] = 1'b1;
      zz_rom_51[4] = 1'b1;
      zz_rom_51[5] = 1'b1;
      zz_rom_51[6] = 1'b1;
      zz_rom_51[7] = 1'b1;
      zz_rom_51[8] = 1'b1;
      zz_rom_51[9] = 1'b1;
      zz_rom_51[10] = 1'b1;
      zz_rom_51[11] = 1'b1;
      zz_rom_51[12] = 1'b1;
      zz_rom_51[13] = 1'b1;
      zz_rom_51[14] = 1'b1;
      zz_rom_51[15] = 1'b1;
      zz_rom_51[16] = 1'b1;
      zz_rom_51[17] = 1'b1;
      zz_rom_51[18] = 1'b1;
      zz_rom_51[19] = 1'b1;
      zz_rom_51[20] = 1'b1;
      zz_rom_51[21] = 1'b1;
      zz_rom_51[22] = 1'b1;
      zz_rom_51[23] = 1'b1;
      zz_rom_51[24] = 1'b1;
      zz_rom_51[25] = 1'b1;
      zz_rom_51[26] = 1'b1;
      zz_rom_51[27] = 1'b1;
      zz_rom_51[28] = 1'b1;
      zz_rom_51[29] = 1'b1;
      zz_rom_51[30] = 1'b1;
      zz_rom_51[31] = 1'b1;
      zz_rom_51[32] = 1'b1;
      zz_rom_51[33] = 1'b1;
      zz_rom_51[34] = 1'b1;
      zz_rom_51[35] = 1'b1;
      zz_rom_51[36] = 1'b1;
      zz_rom_51[37] = 1'b1;
      zz_rom_51[38] = 1'b1;
      zz_rom_51[39] = 1'b1;
      zz_rom_51[40] = 1'b1;
      zz_rom_51[41] = 1'b1;
      zz_rom_51[42] = 1'b1;
      zz_rom_51[43] = 1'b1;
      zz_rom_51[44] = 1'b1;
      zz_rom_51[45] = 1'b1;
      zz_rom_51[46] = 1'b1;
      zz_rom_51[47] = 1'b1;
      zz_rom_51[48] = 1'b1;
      zz_rom_51[49] = 1'b1;
      zz_rom_51[50] = 1'b1;
      zz_rom_51[51] = 1'b1;
      zz_rom_51[52] = 1'b1;
      zz_rom_51[53] = 1'b1;
      zz_rom_51[54] = 1'b1;
      zz_rom_51[55] = 1'b1;
      zz_rom_51[56] = 1'b1;
      zz_rom_51[57] = 1'b1;
      zz_rom_51[58] = 1'b1;
      zz_rom_51[59] = 1'b1;
      zz_rom_51[60] = 1'b1;
      zz_rom_51[61] = 1'b1;
      zz_rom_51[62] = 1'b1;
      zz_rom_51[63] = 1'b1;
      zz_rom_51[64] = 1'b1;
      zz_rom_51[65] = 1'b1;
      zz_rom_51[66] = 1'b1;
      zz_rom_51[67] = 1'b1;
      zz_rom_51[68] = 1'b1;
      zz_rom_51[69] = 1'b1;
      zz_rom_51[70] = 1'b1;
      zz_rom_51[71] = 1'b1;
      zz_rom_51[72] = 1'b1;
      zz_rom_51[73] = 1'b1;
      zz_rom_51[74] = 1'b1;
      zz_rom_51[75] = 1'b1;
      zz_rom_51[76] = 1'b1;
      zz_rom_51[77] = 1'b1;
      zz_rom_51[78] = 1'b1;
      zz_rom_51[79] = 1'b1;
      zz_rom_51[80] = 1'b1;
      zz_rom_51[81] = 1'b1;
      zz_rom_51[82] = 1'b1;
      zz_rom_51[83] = 1'b1;
      zz_rom_51[84] = 1'b1;
      zz_rom_51[85] = 1'b1;
      zz_rom_51[86] = 1'b1;
      zz_rom_51[87] = 1'b1;
      zz_rom_51[88] = 1'b1;
      zz_rom_51[89] = 1'b1;
      zz_rom_51[90] = 1'b1;
      zz_rom_51[91] = 1'b1;
      zz_rom_51[92] = 1'b1;
      zz_rom_51[93] = 1'b1;
      zz_rom_51[94] = 1'b1;
      zz_rom_51[95] = 1'b1;
      zz_rom_51[96] = 1'b1;
      zz_rom_51[97] = 1'b1;
      zz_rom_51[98] = 1'b1;
      zz_rom_51[99] = 1'b1;
    end
  endfunction
  wire [99:0] _zz_52;
  function [99:0] zz_rom_52(input dummy);
    begin
      zz_rom_52[0] = 1'b0;
      zz_rom_52[1] = 1'b1;
      zz_rom_52[2] = 1'b1;
      zz_rom_52[3] = 1'b1;
      zz_rom_52[4] = 1'b1;
      zz_rom_52[5] = 1'b1;
      zz_rom_52[6] = 1'b1;
      zz_rom_52[7] = 1'b1;
      zz_rom_52[8] = 1'b1;
      zz_rom_52[9] = 1'b1;
      zz_rom_52[10] = 1'b1;
      zz_rom_52[11] = 1'b1;
      zz_rom_52[12] = 1'b1;
      zz_rom_52[13] = 1'b1;
      zz_rom_52[14] = 1'b1;
      zz_rom_52[15] = 1'b1;
      zz_rom_52[16] = 1'b1;
      zz_rom_52[17] = 1'b1;
      zz_rom_52[18] = 1'b1;
      zz_rom_52[19] = 1'b1;
      zz_rom_52[20] = 1'b1;
      zz_rom_52[21] = 1'b1;
      zz_rom_52[22] = 1'b1;
      zz_rom_52[23] = 1'b1;
      zz_rom_52[24] = 1'b1;
      zz_rom_52[25] = 1'b1;
      zz_rom_52[26] = 1'b1;
      zz_rom_52[27] = 1'b1;
      zz_rom_52[28] = 1'b1;
      zz_rom_52[29] = 1'b1;
      zz_rom_52[30] = 1'b1;
      zz_rom_52[31] = 1'b1;
      zz_rom_52[32] = 1'b1;
      zz_rom_52[33] = 1'b1;
      zz_rom_52[34] = 1'b1;
      zz_rom_52[35] = 1'b1;
      zz_rom_52[36] = 1'b1;
      zz_rom_52[37] = 1'b1;
      zz_rom_52[38] = 1'b1;
      zz_rom_52[39] = 1'b1;
      zz_rom_52[40] = 1'b1;
      zz_rom_52[41] = 1'b1;
      zz_rom_52[42] = 1'b1;
      zz_rom_52[43] = 1'b1;
      zz_rom_52[44] = 1'b1;
      zz_rom_52[45] = 1'b1;
      zz_rom_52[46] = 1'b1;
      zz_rom_52[47] = 1'b1;
      zz_rom_52[48] = 1'b1;
      zz_rom_52[49] = 1'b1;
      zz_rom_52[50] = 1'b1;
      zz_rom_52[51] = 1'b1;
      zz_rom_52[52] = 1'b1;
      zz_rom_52[53] = 1'b1;
      zz_rom_52[54] = 1'b1;
      zz_rom_52[55] = 1'b1;
      zz_rom_52[56] = 1'b1;
      zz_rom_52[57] = 1'b1;
      zz_rom_52[58] = 1'b1;
      zz_rom_52[59] = 1'b1;
      zz_rom_52[60] = 1'b1;
      zz_rom_52[61] = 1'b1;
      zz_rom_52[62] = 1'b1;
      zz_rom_52[63] = 1'b1;
      zz_rom_52[64] = 1'b1;
      zz_rom_52[65] = 1'b1;
      zz_rom_52[66] = 1'b1;
      zz_rom_52[67] = 1'b1;
      zz_rom_52[68] = 1'b1;
      zz_rom_52[69] = 1'b1;
      zz_rom_52[70] = 1'b1;
      zz_rom_52[71] = 1'b1;
      zz_rom_52[72] = 1'b1;
      zz_rom_52[73] = 1'b1;
      zz_rom_52[74] = 1'b1;
      zz_rom_52[75] = 1'b1;
      zz_rom_52[76] = 1'b1;
      zz_rom_52[77] = 1'b1;
      zz_rom_52[78] = 1'b1;
      zz_rom_52[79] = 1'b1;
      zz_rom_52[80] = 1'b1;
      zz_rom_52[81] = 1'b1;
      zz_rom_52[82] = 1'b1;
      zz_rom_52[83] = 1'b1;
      zz_rom_52[84] = 1'b1;
      zz_rom_52[85] = 1'b1;
      zz_rom_52[86] = 1'b1;
      zz_rom_52[87] = 1'b1;
      zz_rom_52[88] = 1'b1;
      zz_rom_52[89] = 1'b1;
      zz_rom_52[90] = 1'b1;
      zz_rom_52[91] = 1'b1;
      zz_rom_52[92] = 1'b1;
      zz_rom_52[93] = 1'b1;
      zz_rom_52[94] = 1'b1;
      zz_rom_52[95] = 1'b1;
      zz_rom_52[96] = 1'b1;
      zz_rom_52[97] = 1'b1;
      zz_rom_52[98] = 1'b1;
      zz_rom_52[99] = 1'b1;
    end
  endfunction
  wire [99:0] _zz_53;
  function [99:0] zz_rom_53(input dummy);
    begin
      zz_rom_53[0] = 1'b0;
      zz_rom_53[1] = 1'b1;
      zz_rom_53[2] = 1'b1;
      zz_rom_53[3] = 1'b1;
      zz_rom_53[4] = 1'b1;
      zz_rom_53[5] = 1'b1;
      zz_rom_53[6] = 1'b1;
      zz_rom_53[7] = 1'b1;
      zz_rom_53[8] = 1'b1;
      zz_rom_53[9] = 1'b1;
      zz_rom_53[10] = 1'b1;
      zz_rom_53[11] = 1'b1;
      zz_rom_53[12] = 1'b1;
      zz_rom_53[13] = 1'b1;
      zz_rom_53[14] = 1'b1;
      zz_rom_53[15] = 1'b1;
      zz_rom_53[16] = 1'b1;
      zz_rom_53[17] = 1'b1;
      zz_rom_53[18] = 1'b1;
      zz_rom_53[19] = 1'b1;
      zz_rom_53[20] = 1'b1;
      zz_rom_53[21] = 1'b1;
      zz_rom_53[22] = 1'b1;
      zz_rom_53[23] = 1'b1;
      zz_rom_53[24] = 1'b1;
      zz_rom_53[25] = 1'b1;
      zz_rom_53[26] = 1'b1;
      zz_rom_53[27] = 1'b1;
      zz_rom_53[28] = 1'b1;
      zz_rom_53[29] = 1'b1;
      zz_rom_53[30] = 1'b1;
      zz_rom_53[31] = 1'b1;
      zz_rom_53[32] = 1'b1;
      zz_rom_53[33] = 1'b1;
      zz_rom_53[34] = 1'b1;
      zz_rom_53[35] = 1'b1;
      zz_rom_53[36] = 1'b1;
      zz_rom_53[37] = 1'b1;
      zz_rom_53[38] = 1'b1;
      zz_rom_53[39] = 1'b1;
      zz_rom_53[40] = 1'b1;
      zz_rom_53[41] = 1'b1;
      zz_rom_53[42] = 1'b1;
      zz_rom_53[43] = 1'b1;
      zz_rom_53[44] = 1'b1;
      zz_rom_53[45] = 1'b1;
      zz_rom_53[46] = 1'b1;
      zz_rom_53[47] = 1'b1;
      zz_rom_53[48] = 1'b1;
      zz_rom_53[49] = 1'b1;
      zz_rom_53[50] = 1'b1;
      zz_rom_53[51] = 1'b1;
      zz_rom_53[52] = 1'b1;
      zz_rom_53[53] = 1'b1;
      zz_rom_53[54] = 1'b1;
      zz_rom_53[55] = 1'b1;
      zz_rom_53[56] = 1'b1;
      zz_rom_53[57] = 1'b1;
      zz_rom_53[58] = 1'b1;
      zz_rom_53[59] = 1'b1;
      zz_rom_53[60] = 1'b1;
      zz_rom_53[61] = 1'b1;
      zz_rom_53[62] = 1'b1;
      zz_rom_53[63] = 1'b1;
      zz_rom_53[64] = 1'b1;
      zz_rom_53[65] = 1'b1;
      zz_rom_53[66] = 1'b1;
      zz_rom_53[67] = 1'b1;
      zz_rom_53[68] = 1'b1;
      zz_rom_53[69] = 1'b1;
      zz_rom_53[70] = 1'b1;
      zz_rom_53[71] = 1'b1;
      zz_rom_53[72] = 1'b1;
      zz_rom_53[73] = 1'b1;
      zz_rom_53[74] = 1'b1;
      zz_rom_53[75] = 1'b1;
      zz_rom_53[76] = 1'b1;
      zz_rom_53[77] = 1'b1;
      zz_rom_53[78] = 1'b1;
      zz_rom_53[79] = 1'b1;
      zz_rom_53[80] = 1'b1;
      zz_rom_53[81] = 1'b1;
      zz_rom_53[82] = 1'b1;
      zz_rom_53[83] = 1'b1;
      zz_rom_53[84] = 1'b1;
      zz_rom_53[85] = 1'b1;
      zz_rom_53[86] = 1'b1;
      zz_rom_53[87] = 1'b1;
      zz_rom_53[88] = 1'b1;
      zz_rom_53[89] = 1'b1;
      zz_rom_53[90] = 1'b1;
      zz_rom_53[91] = 1'b1;
      zz_rom_53[92] = 1'b1;
      zz_rom_53[93] = 1'b1;
      zz_rom_53[94] = 1'b1;
      zz_rom_53[95] = 1'b1;
      zz_rom_53[96] = 1'b1;
      zz_rom_53[97] = 1'b1;
      zz_rom_53[98] = 1'b1;
      zz_rom_53[99] = 1'b1;
    end
  endfunction
  wire [99:0] _zz_54;
  function [99:0] zz_rom_54(input dummy);
    begin
      zz_rom_54[0] = 1'b0;
      zz_rom_54[1] = 1'b1;
      zz_rom_54[2] = 1'b1;
      zz_rom_54[3] = 1'b1;
      zz_rom_54[4] = 1'b1;
      zz_rom_54[5] = 1'b1;
      zz_rom_54[6] = 1'b1;
      zz_rom_54[7] = 1'b1;
      zz_rom_54[8] = 1'b1;
      zz_rom_54[9] = 1'b1;
      zz_rom_54[10] = 1'b1;
      zz_rom_54[11] = 1'b1;
      zz_rom_54[12] = 1'b1;
      zz_rom_54[13] = 1'b1;
      zz_rom_54[14] = 1'b1;
      zz_rom_54[15] = 1'b1;
      zz_rom_54[16] = 1'b1;
      zz_rom_54[17] = 1'b1;
      zz_rom_54[18] = 1'b1;
      zz_rom_54[19] = 1'b1;
      zz_rom_54[20] = 1'b1;
      zz_rom_54[21] = 1'b1;
      zz_rom_54[22] = 1'b1;
      zz_rom_54[23] = 1'b1;
      zz_rom_54[24] = 1'b1;
      zz_rom_54[25] = 1'b1;
      zz_rom_54[26] = 1'b1;
      zz_rom_54[27] = 1'b1;
      zz_rom_54[28] = 1'b1;
      zz_rom_54[29] = 1'b1;
      zz_rom_54[30] = 1'b1;
      zz_rom_54[31] = 1'b1;
      zz_rom_54[32] = 1'b1;
      zz_rom_54[33] = 1'b1;
      zz_rom_54[34] = 1'b1;
      zz_rom_54[35] = 1'b1;
      zz_rom_54[36] = 1'b1;
      zz_rom_54[37] = 1'b1;
      zz_rom_54[38] = 1'b1;
      zz_rom_54[39] = 1'b1;
      zz_rom_54[40] = 1'b1;
      zz_rom_54[41] = 1'b1;
      zz_rom_54[42] = 1'b1;
      zz_rom_54[43] = 1'b1;
      zz_rom_54[44] = 1'b1;
      zz_rom_54[45] = 1'b1;
      zz_rom_54[46] = 1'b1;
      zz_rom_54[47] = 1'b1;
      zz_rom_54[48] = 1'b1;
      zz_rom_54[49] = 1'b1;
      zz_rom_54[50] = 1'b1;
      zz_rom_54[51] = 1'b1;
      zz_rom_54[52] = 1'b1;
      zz_rom_54[53] = 1'b1;
      zz_rom_54[54] = 1'b1;
      zz_rom_54[55] = 1'b1;
      zz_rom_54[56] = 1'b1;
      zz_rom_54[57] = 1'b1;
      zz_rom_54[58] = 1'b1;
      zz_rom_54[59] = 1'b1;
      zz_rom_54[60] = 1'b1;
      zz_rom_54[61] = 1'b1;
      zz_rom_54[62] = 1'b1;
      zz_rom_54[63] = 1'b1;
      zz_rom_54[64] = 1'b1;
      zz_rom_54[65] = 1'b1;
      zz_rom_54[66] = 1'b1;
      zz_rom_54[67] = 1'b1;
      zz_rom_54[68] = 1'b1;
      zz_rom_54[69] = 1'b1;
      zz_rom_54[70] = 1'b1;
      zz_rom_54[71] = 1'b1;
      zz_rom_54[72] = 1'b1;
      zz_rom_54[73] = 1'b1;
      zz_rom_54[74] = 1'b1;
      zz_rom_54[75] = 1'b1;
      zz_rom_54[76] = 1'b1;
      zz_rom_54[77] = 1'b1;
      zz_rom_54[78] = 1'b1;
      zz_rom_54[79] = 1'b1;
      zz_rom_54[80] = 1'b1;
      zz_rom_54[81] = 1'b1;
      zz_rom_54[82] = 1'b1;
      zz_rom_54[83] = 1'b1;
      zz_rom_54[84] = 1'b1;
      zz_rom_54[85] = 1'b1;
      zz_rom_54[86] = 1'b1;
      zz_rom_54[87] = 1'b1;
      zz_rom_54[88] = 1'b1;
      zz_rom_54[89] = 1'b1;
      zz_rom_54[90] = 1'b1;
      zz_rom_54[91] = 1'b1;
      zz_rom_54[92] = 1'b1;
      zz_rom_54[93] = 1'b1;
      zz_rom_54[94] = 1'b1;
      zz_rom_54[95] = 1'b1;
      zz_rom_54[96] = 1'b1;
      zz_rom_54[97] = 1'b1;
      zz_rom_54[98] = 1'b1;
      zz_rom_54[99] = 1'b1;
    end
  endfunction
  wire [99:0] _zz_55;
  function [99:0] zz_rom_55(input dummy);
    begin
      zz_rom_55[0] = 1'b0;
      zz_rom_55[1] = 1'b1;
      zz_rom_55[2] = 1'b1;
      zz_rom_55[3] = 1'b1;
      zz_rom_55[4] = 1'b1;
      zz_rom_55[5] = 1'b1;
      zz_rom_55[6] = 1'b1;
      zz_rom_55[7] = 1'b1;
      zz_rom_55[8] = 1'b1;
      zz_rom_55[9] = 1'b1;
      zz_rom_55[10] = 1'b1;
      zz_rom_55[11] = 1'b1;
      zz_rom_55[12] = 1'b1;
      zz_rom_55[13] = 1'b1;
      zz_rom_55[14] = 1'b1;
      zz_rom_55[15] = 1'b1;
      zz_rom_55[16] = 1'b1;
      zz_rom_55[17] = 1'b1;
      zz_rom_55[18] = 1'b1;
      zz_rom_55[19] = 1'b1;
      zz_rom_55[20] = 1'b1;
      zz_rom_55[21] = 1'b1;
      zz_rom_55[22] = 1'b1;
      zz_rom_55[23] = 1'b1;
      zz_rom_55[24] = 1'b1;
      zz_rom_55[25] = 1'b1;
      zz_rom_55[26] = 1'b1;
      zz_rom_55[27] = 1'b1;
      zz_rom_55[28] = 1'b1;
      zz_rom_55[29] = 1'b1;
      zz_rom_55[30] = 1'b1;
      zz_rom_55[31] = 1'b1;
      zz_rom_55[32] = 1'b1;
      zz_rom_55[33] = 1'b1;
      zz_rom_55[34] = 1'b1;
      zz_rom_55[35] = 1'b1;
      zz_rom_55[36] = 1'b1;
      zz_rom_55[37] = 1'b1;
      zz_rom_55[38] = 1'b1;
      zz_rom_55[39] = 1'b1;
      zz_rom_55[40] = 1'b1;
      zz_rom_55[41] = 1'b1;
      zz_rom_55[42] = 1'b1;
      zz_rom_55[43] = 1'b1;
      zz_rom_55[44] = 1'b1;
      zz_rom_55[45] = 1'b1;
      zz_rom_55[46] = 1'b1;
      zz_rom_55[47] = 1'b1;
      zz_rom_55[48] = 1'b1;
      zz_rom_55[49] = 1'b1;
      zz_rom_55[50] = 1'b1;
      zz_rom_55[51] = 1'b1;
      zz_rom_55[52] = 1'b1;
      zz_rom_55[53] = 1'b1;
      zz_rom_55[54] = 1'b1;
      zz_rom_55[55] = 1'b1;
      zz_rom_55[56] = 1'b1;
      zz_rom_55[57] = 1'b1;
      zz_rom_55[58] = 1'b1;
      zz_rom_55[59] = 1'b1;
      zz_rom_55[60] = 1'b1;
      zz_rom_55[61] = 1'b1;
      zz_rom_55[62] = 1'b1;
      zz_rom_55[63] = 1'b1;
      zz_rom_55[64] = 1'b1;
      zz_rom_55[65] = 1'b1;
      zz_rom_55[66] = 1'b1;
      zz_rom_55[67] = 1'b1;
      zz_rom_55[68] = 1'b1;
      zz_rom_55[69] = 1'b1;
      zz_rom_55[70] = 1'b1;
      zz_rom_55[71] = 1'b1;
      zz_rom_55[72] = 1'b1;
      zz_rom_55[73] = 1'b1;
      zz_rom_55[74] = 1'b1;
      zz_rom_55[75] = 1'b1;
      zz_rom_55[76] = 1'b1;
      zz_rom_55[77] = 1'b1;
      zz_rom_55[78] = 1'b1;
      zz_rom_55[79] = 1'b1;
      zz_rom_55[80] = 1'b1;
      zz_rom_55[81] = 1'b1;
      zz_rom_55[82] = 1'b1;
      zz_rom_55[83] = 1'b1;
      zz_rom_55[84] = 1'b1;
      zz_rom_55[85] = 1'b1;
      zz_rom_55[86] = 1'b1;
      zz_rom_55[87] = 1'b1;
      zz_rom_55[88] = 1'b1;
      zz_rom_55[89] = 1'b1;
      zz_rom_55[90] = 1'b1;
      zz_rom_55[91] = 1'b1;
      zz_rom_55[92] = 1'b1;
      zz_rom_55[93] = 1'b1;
      zz_rom_55[94] = 1'b1;
      zz_rom_55[95] = 1'b1;
      zz_rom_55[96] = 1'b1;
      zz_rom_55[97] = 1'b1;
      zz_rom_55[98] = 1'b1;
      zz_rom_55[99] = 1'b1;
    end
  endfunction
  wire [99:0] _zz_56;
  function [99:0] zz_rom_56(input dummy);
    begin
      zz_rom_56[0] = 1'b0;
      zz_rom_56[1] = 1'b1;
      zz_rom_56[2] = 1'b1;
      zz_rom_56[3] = 1'b1;
      zz_rom_56[4] = 1'b1;
      zz_rom_56[5] = 1'b1;
      zz_rom_56[6] = 1'b1;
      zz_rom_56[7] = 1'b1;
      zz_rom_56[8] = 1'b1;
      zz_rom_56[9] = 1'b1;
      zz_rom_56[10] = 1'b1;
      zz_rom_56[11] = 1'b1;
      zz_rom_56[12] = 1'b1;
      zz_rom_56[13] = 1'b1;
      zz_rom_56[14] = 1'b1;
      zz_rom_56[15] = 1'b1;
      zz_rom_56[16] = 1'b1;
      zz_rom_56[17] = 1'b1;
      zz_rom_56[18] = 1'b1;
      zz_rom_56[19] = 1'b1;
      zz_rom_56[20] = 1'b1;
      zz_rom_56[21] = 1'b1;
      zz_rom_56[22] = 1'b1;
      zz_rom_56[23] = 1'b1;
      zz_rom_56[24] = 1'b1;
      zz_rom_56[25] = 1'b1;
      zz_rom_56[26] = 1'b1;
      zz_rom_56[27] = 1'b1;
      zz_rom_56[28] = 1'b1;
      zz_rom_56[29] = 1'b1;
      zz_rom_56[30] = 1'b1;
      zz_rom_56[31] = 1'b1;
      zz_rom_56[32] = 1'b1;
      zz_rom_56[33] = 1'b1;
      zz_rom_56[34] = 1'b1;
      zz_rom_56[35] = 1'b1;
      zz_rom_56[36] = 1'b1;
      zz_rom_56[37] = 1'b1;
      zz_rom_56[38] = 1'b1;
      zz_rom_56[39] = 1'b1;
      zz_rom_56[40] = 1'b1;
      zz_rom_56[41] = 1'b1;
      zz_rom_56[42] = 1'b1;
      zz_rom_56[43] = 1'b1;
      zz_rom_56[44] = 1'b1;
      zz_rom_56[45] = 1'b1;
      zz_rom_56[46] = 1'b1;
      zz_rom_56[47] = 1'b1;
      zz_rom_56[48] = 1'b1;
      zz_rom_56[49] = 1'b1;
      zz_rom_56[50] = 1'b1;
      zz_rom_56[51] = 1'b1;
      zz_rom_56[52] = 1'b1;
      zz_rom_56[53] = 1'b1;
      zz_rom_56[54] = 1'b1;
      zz_rom_56[55] = 1'b1;
      zz_rom_56[56] = 1'b1;
      zz_rom_56[57] = 1'b1;
      zz_rom_56[58] = 1'b1;
      zz_rom_56[59] = 1'b1;
      zz_rom_56[60] = 1'b1;
      zz_rom_56[61] = 1'b1;
      zz_rom_56[62] = 1'b1;
      zz_rom_56[63] = 1'b1;
      zz_rom_56[64] = 1'b1;
      zz_rom_56[65] = 1'b1;
      zz_rom_56[66] = 1'b1;
      zz_rom_56[67] = 1'b1;
      zz_rom_56[68] = 1'b1;
      zz_rom_56[69] = 1'b1;
      zz_rom_56[70] = 1'b1;
      zz_rom_56[71] = 1'b1;
      zz_rom_56[72] = 1'b1;
      zz_rom_56[73] = 1'b1;
      zz_rom_56[74] = 1'b1;
      zz_rom_56[75] = 1'b1;
      zz_rom_56[76] = 1'b1;
      zz_rom_56[77] = 1'b1;
      zz_rom_56[78] = 1'b1;
      zz_rom_56[79] = 1'b1;
      zz_rom_56[80] = 1'b1;
      zz_rom_56[81] = 1'b1;
      zz_rom_56[82] = 1'b1;
      zz_rom_56[83] = 1'b1;
      zz_rom_56[84] = 1'b1;
      zz_rom_56[85] = 1'b1;
      zz_rom_56[86] = 1'b1;
      zz_rom_56[87] = 1'b1;
      zz_rom_56[88] = 1'b1;
      zz_rom_56[89] = 1'b1;
      zz_rom_56[90] = 1'b1;
      zz_rom_56[91] = 1'b1;
      zz_rom_56[92] = 1'b1;
      zz_rom_56[93] = 1'b1;
      zz_rom_56[94] = 1'b1;
      zz_rom_56[95] = 1'b1;
      zz_rom_56[96] = 1'b1;
      zz_rom_56[97] = 1'b1;
      zz_rom_56[98] = 1'b1;
      zz_rom_56[99] = 1'b1;
    end
  endfunction
  wire [99:0] _zz_57;
  function [99:0] zz_rom_57(input dummy);
    begin
      zz_rom_57[0] = 1'b0;
      zz_rom_57[1] = 1'b1;
      zz_rom_57[2] = 1'b1;
      zz_rom_57[3] = 1'b1;
      zz_rom_57[4] = 1'b1;
      zz_rom_57[5] = 1'b1;
      zz_rom_57[6] = 1'b1;
      zz_rom_57[7] = 1'b1;
      zz_rom_57[8] = 1'b1;
      zz_rom_57[9] = 1'b1;
      zz_rom_57[10] = 1'b1;
      zz_rom_57[11] = 1'b1;
      zz_rom_57[12] = 1'b1;
      zz_rom_57[13] = 1'b1;
      zz_rom_57[14] = 1'b1;
      zz_rom_57[15] = 1'b1;
      zz_rom_57[16] = 1'b1;
      zz_rom_57[17] = 1'b1;
      zz_rom_57[18] = 1'b1;
      zz_rom_57[19] = 1'b1;
      zz_rom_57[20] = 1'b1;
      zz_rom_57[21] = 1'b1;
      zz_rom_57[22] = 1'b1;
      zz_rom_57[23] = 1'b1;
      zz_rom_57[24] = 1'b1;
      zz_rom_57[25] = 1'b1;
      zz_rom_57[26] = 1'b1;
      zz_rom_57[27] = 1'b1;
      zz_rom_57[28] = 1'b1;
      zz_rom_57[29] = 1'b1;
      zz_rom_57[30] = 1'b1;
      zz_rom_57[31] = 1'b1;
      zz_rom_57[32] = 1'b1;
      zz_rom_57[33] = 1'b1;
      zz_rom_57[34] = 1'b1;
      zz_rom_57[35] = 1'b1;
      zz_rom_57[36] = 1'b1;
      zz_rom_57[37] = 1'b1;
      zz_rom_57[38] = 1'b1;
      zz_rom_57[39] = 1'b1;
      zz_rom_57[40] = 1'b1;
      zz_rom_57[41] = 1'b1;
      zz_rom_57[42] = 1'b1;
      zz_rom_57[43] = 1'b1;
      zz_rom_57[44] = 1'b1;
      zz_rom_57[45] = 1'b1;
      zz_rom_57[46] = 1'b1;
      zz_rom_57[47] = 1'b1;
      zz_rom_57[48] = 1'b1;
      zz_rom_57[49] = 1'b1;
      zz_rom_57[50] = 1'b1;
      zz_rom_57[51] = 1'b1;
      zz_rom_57[52] = 1'b1;
      zz_rom_57[53] = 1'b1;
      zz_rom_57[54] = 1'b1;
      zz_rom_57[55] = 1'b1;
      zz_rom_57[56] = 1'b1;
      zz_rom_57[57] = 1'b1;
      zz_rom_57[58] = 1'b1;
      zz_rom_57[59] = 1'b1;
      zz_rom_57[60] = 1'b1;
      zz_rom_57[61] = 1'b1;
      zz_rom_57[62] = 1'b1;
      zz_rom_57[63] = 1'b1;
      zz_rom_57[64] = 1'b1;
      zz_rom_57[65] = 1'b1;
      zz_rom_57[66] = 1'b1;
      zz_rom_57[67] = 1'b1;
      zz_rom_57[68] = 1'b1;
      zz_rom_57[69] = 1'b1;
      zz_rom_57[70] = 1'b1;
      zz_rom_57[71] = 1'b1;
      zz_rom_57[72] = 1'b1;
      zz_rom_57[73] = 1'b1;
      zz_rom_57[74] = 1'b1;
      zz_rom_57[75] = 1'b1;
      zz_rom_57[76] = 1'b1;
      zz_rom_57[77] = 1'b1;
      zz_rom_57[78] = 1'b1;
      zz_rom_57[79] = 1'b1;
      zz_rom_57[80] = 1'b1;
      zz_rom_57[81] = 1'b1;
      zz_rom_57[82] = 1'b1;
      zz_rom_57[83] = 1'b1;
      zz_rom_57[84] = 1'b1;
      zz_rom_57[85] = 1'b1;
      zz_rom_57[86] = 1'b1;
      zz_rom_57[87] = 1'b1;
      zz_rom_57[88] = 1'b1;
      zz_rom_57[89] = 1'b1;
      zz_rom_57[90] = 1'b1;
      zz_rom_57[91] = 1'b1;
      zz_rom_57[92] = 1'b1;
      zz_rom_57[93] = 1'b1;
      zz_rom_57[94] = 1'b1;
      zz_rom_57[95] = 1'b1;
      zz_rom_57[96] = 1'b1;
      zz_rom_57[97] = 1'b1;
      zz_rom_57[98] = 1'b1;
      zz_rom_57[99] = 1'b1;
    end
  endfunction
  wire [99:0] _zz_58;
  function [99:0] zz_rom_58(input dummy);
    begin
      zz_rom_58[0] = 1'b0;
      zz_rom_58[1] = 1'b1;
      zz_rom_58[2] = 1'b1;
      zz_rom_58[3] = 1'b1;
      zz_rom_58[4] = 1'b1;
      zz_rom_58[5] = 1'b1;
      zz_rom_58[6] = 1'b1;
      zz_rom_58[7] = 1'b1;
      zz_rom_58[8] = 1'b1;
      zz_rom_58[9] = 1'b1;
      zz_rom_58[10] = 1'b1;
      zz_rom_58[11] = 1'b1;
      zz_rom_58[12] = 1'b1;
      zz_rom_58[13] = 1'b1;
      zz_rom_58[14] = 1'b1;
      zz_rom_58[15] = 1'b1;
      zz_rom_58[16] = 1'b1;
      zz_rom_58[17] = 1'b1;
      zz_rom_58[18] = 1'b1;
      zz_rom_58[19] = 1'b1;
      zz_rom_58[20] = 1'b1;
      zz_rom_58[21] = 1'b1;
      zz_rom_58[22] = 1'b1;
      zz_rom_58[23] = 1'b1;
      zz_rom_58[24] = 1'b1;
      zz_rom_58[25] = 1'b1;
      zz_rom_58[26] = 1'b1;
      zz_rom_58[27] = 1'b1;
      zz_rom_58[28] = 1'b1;
      zz_rom_58[29] = 1'b1;
      zz_rom_58[30] = 1'b1;
      zz_rom_58[31] = 1'b1;
      zz_rom_58[32] = 1'b1;
      zz_rom_58[33] = 1'b1;
      zz_rom_58[34] = 1'b1;
      zz_rom_58[35] = 1'b1;
      zz_rom_58[36] = 1'b1;
      zz_rom_58[37] = 1'b1;
      zz_rom_58[38] = 1'b1;
      zz_rom_58[39] = 1'b1;
      zz_rom_58[40] = 1'b1;
      zz_rom_58[41] = 1'b1;
      zz_rom_58[42] = 1'b1;
      zz_rom_58[43] = 1'b1;
      zz_rom_58[44] = 1'b1;
      zz_rom_58[45] = 1'b1;
      zz_rom_58[46] = 1'b1;
      zz_rom_58[47] = 1'b1;
      zz_rom_58[48] = 1'b1;
      zz_rom_58[49] = 1'b1;
      zz_rom_58[50] = 1'b1;
      zz_rom_58[51] = 1'b1;
      zz_rom_58[52] = 1'b1;
      zz_rom_58[53] = 1'b1;
      zz_rom_58[54] = 1'b1;
      zz_rom_58[55] = 1'b1;
      zz_rom_58[56] = 1'b1;
      zz_rom_58[57] = 1'b1;
      zz_rom_58[58] = 1'b1;
      zz_rom_58[59] = 1'b1;
      zz_rom_58[60] = 1'b1;
      zz_rom_58[61] = 1'b1;
      zz_rom_58[62] = 1'b1;
      zz_rom_58[63] = 1'b1;
      zz_rom_58[64] = 1'b1;
      zz_rom_58[65] = 1'b1;
      zz_rom_58[66] = 1'b1;
      zz_rom_58[67] = 1'b1;
      zz_rom_58[68] = 1'b1;
      zz_rom_58[69] = 1'b1;
      zz_rom_58[70] = 1'b1;
      zz_rom_58[71] = 1'b1;
      zz_rom_58[72] = 1'b1;
      zz_rom_58[73] = 1'b1;
      zz_rom_58[74] = 1'b1;
      zz_rom_58[75] = 1'b1;
      zz_rom_58[76] = 1'b1;
      zz_rom_58[77] = 1'b1;
      zz_rom_58[78] = 1'b1;
      zz_rom_58[79] = 1'b1;
      zz_rom_58[80] = 1'b1;
      zz_rom_58[81] = 1'b1;
      zz_rom_58[82] = 1'b1;
      zz_rom_58[83] = 1'b1;
      zz_rom_58[84] = 1'b1;
      zz_rom_58[85] = 1'b1;
      zz_rom_58[86] = 1'b1;
      zz_rom_58[87] = 1'b1;
      zz_rom_58[88] = 1'b1;
      zz_rom_58[89] = 1'b1;
      zz_rom_58[90] = 1'b1;
      zz_rom_58[91] = 1'b1;
      zz_rom_58[92] = 1'b1;
      zz_rom_58[93] = 1'b1;
      zz_rom_58[94] = 1'b1;
      zz_rom_58[95] = 1'b1;
      zz_rom_58[96] = 1'b1;
      zz_rom_58[97] = 1'b1;
      zz_rom_58[98] = 1'b1;
      zz_rom_58[99] = 1'b1;
    end
  endfunction
  wire [99:0] _zz_59;
  function [99:0] zz_rom_59(input dummy);
    begin
      zz_rom_59[0] = 1'b0;
      zz_rom_59[1] = 1'b1;
      zz_rom_59[2] = 1'b1;
      zz_rom_59[3] = 1'b1;
      zz_rom_59[4] = 1'b1;
      zz_rom_59[5] = 1'b1;
      zz_rom_59[6] = 1'b1;
      zz_rom_59[7] = 1'b1;
      zz_rom_59[8] = 1'b1;
      zz_rom_59[9] = 1'b1;
      zz_rom_59[10] = 1'b1;
      zz_rom_59[11] = 1'b1;
      zz_rom_59[12] = 1'b1;
      zz_rom_59[13] = 1'b1;
      zz_rom_59[14] = 1'b1;
      zz_rom_59[15] = 1'b1;
      zz_rom_59[16] = 1'b1;
      zz_rom_59[17] = 1'b1;
      zz_rom_59[18] = 1'b1;
      zz_rom_59[19] = 1'b1;
      zz_rom_59[20] = 1'b1;
      zz_rom_59[21] = 1'b1;
      zz_rom_59[22] = 1'b1;
      zz_rom_59[23] = 1'b1;
      zz_rom_59[24] = 1'b1;
      zz_rom_59[25] = 1'b1;
      zz_rom_59[26] = 1'b1;
      zz_rom_59[27] = 1'b1;
      zz_rom_59[28] = 1'b1;
      zz_rom_59[29] = 1'b1;
      zz_rom_59[30] = 1'b1;
      zz_rom_59[31] = 1'b1;
      zz_rom_59[32] = 1'b1;
      zz_rom_59[33] = 1'b1;
      zz_rom_59[34] = 1'b1;
      zz_rom_59[35] = 1'b1;
      zz_rom_59[36] = 1'b1;
      zz_rom_59[37] = 1'b1;
      zz_rom_59[38] = 1'b1;
      zz_rom_59[39] = 1'b1;
      zz_rom_59[40] = 1'b1;
      zz_rom_59[41] = 1'b1;
      zz_rom_59[42] = 1'b1;
      zz_rom_59[43] = 1'b1;
      zz_rom_59[44] = 1'b1;
      zz_rom_59[45] = 1'b1;
      zz_rom_59[46] = 1'b1;
      zz_rom_59[47] = 1'b1;
      zz_rom_59[48] = 1'b1;
      zz_rom_59[49] = 1'b1;
      zz_rom_59[50] = 1'b1;
      zz_rom_59[51] = 1'b1;
      zz_rom_59[52] = 1'b1;
      zz_rom_59[53] = 1'b1;
      zz_rom_59[54] = 1'b1;
      zz_rom_59[55] = 1'b1;
      zz_rom_59[56] = 1'b1;
      zz_rom_59[57] = 1'b1;
      zz_rom_59[58] = 1'b1;
      zz_rom_59[59] = 1'b1;
      zz_rom_59[60] = 1'b1;
      zz_rom_59[61] = 1'b1;
      zz_rom_59[62] = 1'b1;
      zz_rom_59[63] = 1'b1;
      zz_rom_59[64] = 1'b1;
      zz_rom_59[65] = 1'b1;
      zz_rom_59[66] = 1'b1;
      zz_rom_59[67] = 1'b1;
      zz_rom_59[68] = 1'b1;
      zz_rom_59[69] = 1'b1;
      zz_rom_59[70] = 1'b1;
      zz_rom_59[71] = 1'b1;
      zz_rom_59[72] = 1'b1;
      zz_rom_59[73] = 1'b1;
      zz_rom_59[74] = 1'b1;
      zz_rom_59[75] = 1'b1;
      zz_rom_59[76] = 1'b1;
      zz_rom_59[77] = 1'b1;
      zz_rom_59[78] = 1'b1;
      zz_rom_59[79] = 1'b1;
      zz_rom_59[80] = 1'b1;
      zz_rom_59[81] = 1'b1;
      zz_rom_59[82] = 1'b1;
      zz_rom_59[83] = 1'b1;
      zz_rom_59[84] = 1'b1;
      zz_rom_59[85] = 1'b1;
      zz_rom_59[86] = 1'b1;
      zz_rom_59[87] = 1'b1;
      zz_rom_59[88] = 1'b1;
      zz_rom_59[89] = 1'b1;
      zz_rom_59[90] = 1'b1;
      zz_rom_59[91] = 1'b1;
      zz_rom_59[92] = 1'b1;
      zz_rom_59[93] = 1'b1;
      zz_rom_59[94] = 1'b1;
      zz_rom_59[95] = 1'b1;
      zz_rom_59[96] = 1'b1;
      zz_rom_59[97] = 1'b1;
      zz_rom_59[98] = 1'b1;
      zz_rom_59[99] = 1'b1;
    end
  endfunction
  wire [99:0] _zz_60;
  function [99:0] zz_rom_60(input dummy);
    begin
      zz_rom_60[0] = 1'b0;
      zz_rom_60[1] = 1'b0;
      zz_rom_60[2] = 1'b1;
      zz_rom_60[3] = 1'b1;
      zz_rom_60[4] = 1'b1;
      zz_rom_60[5] = 1'b1;
      zz_rom_60[6] = 1'b1;
      zz_rom_60[7] = 1'b1;
      zz_rom_60[8] = 1'b1;
      zz_rom_60[9] = 1'b1;
      zz_rom_60[10] = 1'b1;
      zz_rom_60[11] = 1'b1;
      zz_rom_60[12] = 1'b1;
      zz_rom_60[13] = 1'b1;
      zz_rom_60[14] = 1'b1;
      zz_rom_60[15] = 1'b1;
      zz_rom_60[16] = 1'b1;
      zz_rom_60[17] = 1'b1;
      zz_rom_60[18] = 1'b1;
      zz_rom_60[19] = 1'b1;
      zz_rom_60[20] = 1'b1;
      zz_rom_60[21] = 1'b1;
      zz_rom_60[22] = 1'b1;
      zz_rom_60[23] = 1'b1;
      zz_rom_60[24] = 1'b1;
      zz_rom_60[25] = 1'b1;
      zz_rom_60[26] = 1'b1;
      zz_rom_60[27] = 1'b1;
      zz_rom_60[28] = 1'b1;
      zz_rom_60[29] = 1'b1;
      zz_rom_60[30] = 1'b1;
      zz_rom_60[31] = 1'b1;
      zz_rom_60[32] = 1'b1;
      zz_rom_60[33] = 1'b1;
      zz_rom_60[34] = 1'b1;
      zz_rom_60[35] = 1'b1;
      zz_rom_60[36] = 1'b1;
      zz_rom_60[37] = 1'b1;
      zz_rom_60[38] = 1'b1;
      zz_rom_60[39] = 1'b1;
      zz_rom_60[40] = 1'b1;
      zz_rom_60[41] = 1'b1;
      zz_rom_60[42] = 1'b1;
      zz_rom_60[43] = 1'b1;
      zz_rom_60[44] = 1'b1;
      zz_rom_60[45] = 1'b1;
      zz_rom_60[46] = 1'b1;
      zz_rom_60[47] = 1'b1;
      zz_rom_60[48] = 1'b1;
      zz_rom_60[49] = 1'b1;
      zz_rom_60[50] = 1'b1;
      zz_rom_60[51] = 1'b1;
      zz_rom_60[52] = 1'b1;
      zz_rom_60[53] = 1'b1;
      zz_rom_60[54] = 1'b1;
      zz_rom_60[55] = 1'b1;
      zz_rom_60[56] = 1'b1;
      zz_rom_60[57] = 1'b1;
      zz_rom_60[58] = 1'b1;
      zz_rom_60[59] = 1'b1;
      zz_rom_60[60] = 1'b1;
      zz_rom_60[61] = 1'b1;
      zz_rom_60[62] = 1'b1;
      zz_rom_60[63] = 1'b1;
      zz_rom_60[64] = 1'b1;
      zz_rom_60[65] = 1'b1;
      zz_rom_60[66] = 1'b1;
      zz_rom_60[67] = 1'b1;
      zz_rom_60[68] = 1'b1;
      zz_rom_60[69] = 1'b1;
      zz_rom_60[70] = 1'b1;
      zz_rom_60[71] = 1'b1;
      zz_rom_60[72] = 1'b1;
      zz_rom_60[73] = 1'b1;
      zz_rom_60[74] = 1'b1;
      zz_rom_60[75] = 1'b1;
      zz_rom_60[76] = 1'b1;
      zz_rom_60[77] = 1'b1;
      zz_rom_60[78] = 1'b1;
      zz_rom_60[79] = 1'b1;
      zz_rom_60[80] = 1'b1;
      zz_rom_60[81] = 1'b1;
      zz_rom_60[82] = 1'b1;
      zz_rom_60[83] = 1'b1;
      zz_rom_60[84] = 1'b1;
      zz_rom_60[85] = 1'b1;
      zz_rom_60[86] = 1'b1;
      zz_rom_60[87] = 1'b1;
      zz_rom_60[88] = 1'b1;
      zz_rom_60[89] = 1'b1;
      zz_rom_60[90] = 1'b1;
      zz_rom_60[91] = 1'b1;
      zz_rom_60[92] = 1'b1;
      zz_rom_60[93] = 1'b1;
      zz_rom_60[94] = 1'b1;
      zz_rom_60[95] = 1'b1;
      zz_rom_60[96] = 1'b1;
      zz_rom_60[97] = 1'b1;
      zz_rom_60[98] = 1'b1;
      zz_rom_60[99] = 1'b0;
    end
  endfunction
  wire [99:0] _zz_61;
  function [99:0] zz_rom_61(input dummy);
    begin
      zz_rom_61[0] = 1'b0;
      zz_rom_61[1] = 1'b0;
      zz_rom_61[2] = 1'b1;
      zz_rom_61[3] = 1'b1;
      zz_rom_61[4] = 1'b1;
      zz_rom_61[5] = 1'b1;
      zz_rom_61[6] = 1'b1;
      zz_rom_61[7] = 1'b1;
      zz_rom_61[8] = 1'b1;
      zz_rom_61[9] = 1'b1;
      zz_rom_61[10] = 1'b1;
      zz_rom_61[11] = 1'b1;
      zz_rom_61[12] = 1'b1;
      zz_rom_61[13] = 1'b1;
      zz_rom_61[14] = 1'b1;
      zz_rom_61[15] = 1'b1;
      zz_rom_61[16] = 1'b1;
      zz_rom_61[17] = 1'b1;
      zz_rom_61[18] = 1'b1;
      zz_rom_61[19] = 1'b1;
      zz_rom_61[20] = 1'b1;
      zz_rom_61[21] = 1'b1;
      zz_rom_61[22] = 1'b1;
      zz_rom_61[23] = 1'b1;
      zz_rom_61[24] = 1'b1;
      zz_rom_61[25] = 1'b1;
      zz_rom_61[26] = 1'b1;
      zz_rom_61[27] = 1'b1;
      zz_rom_61[28] = 1'b1;
      zz_rom_61[29] = 1'b1;
      zz_rom_61[30] = 1'b1;
      zz_rom_61[31] = 1'b1;
      zz_rom_61[32] = 1'b1;
      zz_rom_61[33] = 1'b1;
      zz_rom_61[34] = 1'b1;
      zz_rom_61[35] = 1'b1;
      zz_rom_61[36] = 1'b1;
      zz_rom_61[37] = 1'b1;
      zz_rom_61[38] = 1'b1;
      zz_rom_61[39] = 1'b1;
      zz_rom_61[40] = 1'b1;
      zz_rom_61[41] = 1'b1;
      zz_rom_61[42] = 1'b1;
      zz_rom_61[43] = 1'b1;
      zz_rom_61[44] = 1'b1;
      zz_rom_61[45] = 1'b1;
      zz_rom_61[46] = 1'b1;
      zz_rom_61[47] = 1'b1;
      zz_rom_61[48] = 1'b1;
      zz_rom_61[49] = 1'b1;
      zz_rom_61[50] = 1'b1;
      zz_rom_61[51] = 1'b1;
      zz_rom_61[52] = 1'b1;
      zz_rom_61[53] = 1'b1;
      zz_rom_61[54] = 1'b1;
      zz_rom_61[55] = 1'b1;
      zz_rom_61[56] = 1'b1;
      zz_rom_61[57] = 1'b1;
      zz_rom_61[58] = 1'b1;
      zz_rom_61[59] = 1'b1;
      zz_rom_61[60] = 1'b1;
      zz_rom_61[61] = 1'b1;
      zz_rom_61[62] = 1'b1;
      zz_rom_61[63] = 1'b1;
      zz_rom_61[64] = 1'b1;
      zz_rom_61[65] = 1'b1;
      zz_rom_61[66] = 1'b1;
      zz_rom_61[67] = 1'b1;
      zz_rom_61[68] = 1'b1;
      zz_rom_61[69] = 1'b1;
      zz_rom_61[70] = 1'b1;
      zz_rom_61[71] = 1'b1;
      zz_rom_61[72] = 1'b1;
      zz_rom_61[73] = 1'b1;
      zz_rom_61[74] = 1'b1;
      zz_rom_61[75] = 1'b1;
      zz_rom_61[76] = 1'b1;
      zz_rom_61[77] = 1'b1;
      zz_rom_61[78] = 1'b1;
      zz_rom_61[79] = 1'b1;
      zz_rom_61[80] = 1'b1;
      zz_rom_61[81] = 1'b1;
      zz_rom_61[82] = 1'b1;
      zz_rom_61[83] = 1'b1;
      zz_rom_61[84] = 1'b1;
      zz_rom_61[85] = 1'b1;
      zz_rom_61[86] = 1'b1;
      zz_rom_61[87] = 1'b1;
      zz_rom_61[88] = 1'b1;
      zz_rom_61[89] = 1'b1;
      zz_rom_61[90] = 1'b1;
      zz_rom_61[91] = 1'b1;
      zz_rom_61[92] = 1'b1;
      zz_rom_61[93] = 1'b1;
      zz_rom_61[94] = 1'b1;
      zz_rom_61[95] = 1'b1;
      zz_rom_61[96] = 1'b1;
      zz_rom_61[97] = 1'b1;
      zz_rom_61[98] = 1'b1;
      zz_rom_61[99] = 1'b0;
    end
  endfunction
  wire [99:0] _zz_62;
  function [99:0] zz_rom_62(input dummy);
    begin
      zz_rom_62[0] = 1'b0;
      zz_rom_62[1] = 1'b0;
      zz_rom_62[2] = 1'b1;
      zz_rom_62[3] = 1'b1;
      zz_rom_62[4] = 1'b1;
      zz_rom_62[5] = 1'b1;
      zz_rom_62[6] = 1'b1;
      zz_rom_62[7] = 1'b1;
      zz_rom_62[8] = 1'b1;
      zz_rom_62[9] = 1'b1;
      zz_rom_62[10] = 1'b1;
      zz_rom_62[11] = 1'b1;
      zz_rom_62[12] = 1'b1;
      zz_rom_62[13] = 1'b1;
      zz_rom_62[14] = 1'b1;
      zz_rom_62[15] = 1'b1;
      zz_rom_62[16] = 1'b1;
      zz_rom_62[17] = 1'b1;
      zz_rom_62[18] = 1'b1;
      zz_rom_62[19] = 1'b1;
      zz_rom_62[20] = 1'b1;
      zz_rom_62[21] = 1'b1;
      zz_rom_62[22] = 1'b1;
      zz_rom_62[23] = 1'b1;
      zz_rom_62[24] = 1'b1;
      zz_rom_62[25] = 1'b1;
      zz_rom_62[26] = 1'b1;
      zz_rom_62[27] = 1'b1;
      zz_rom_62[28] = 1'b1;
      zz_rom_62[29] = 1'b1;
      zz_rom_62[30] = 1'b1;
      zz_rom_62[31] = 1'b1;
      zz_rom_62[32] = 1'b1;
      zz_rom_62[33] = 1'b1;
      zz_rom_62[34] = 1'b1;
      zz_rom_62[35] = 1'b1;
      zz_rom_62[36] = 1'b1;
      zz_rom_62[37] = 1'b1;
      zz_rom_62[38] = 1'b1;
      zz_rom_62[39] = 1'b1;
      zz_rom_62[40] = 1'b1;
      zz_rom_62[41] = 1'b1;
      zz_rom_62[42] = 1'b1;
      zz_rom_62[43] = 1'b1;
      zz_rom_62[44] = 1'b1;
      zz_rom_62[45] = 1'b1;
      zz_rom_62[46] = 1'b1;
      zz_rom_62[47] = 1'b1;
      zz_rom_62[48] = 1'b1;
      zz_rom_62[49] = 1'b1;
      zz_rom_62[50] = 1'b1;
      zz_rom_62[51] = 1'b1;
      zz_rom_62[52] = 1'b1;
      zz_rom_62[53] = 1'b1;
      zz_rom_62[54] = 1'b1;
      zz_rom_62[55] = 1'b1;
      zz_rom_62[56] = 1'b1;
      zz_rom_62[57] = 1'b1;
      zz_rom_62[58] = 1'b1;
      zz_rom_62[59] = 1'b1;
      zz_rom_62[60] = 1'b1;
      zz_rom_62[61] = 1'b1;
      zz_rom_62[62] = 1'b1;
      zz_rom_62[63] = 1'b1;
      zz_rom_62[64] = 1'b1;
      zz_rom_62[65] = 1'b1;
      zz_rom_62[66] = 1'b1;
      zz_rom_62[67] = 1'b1;
      zz_rom_62[68] = 1'b1;
      zz_rom_62[69] = 1'b1;
      zz_rom_62[70] = 1'b1;
      zz_rom_62[71] = 1'b1;
      zz_rom_62[72] = 1'b1;
      zz_rom_62[73] = 1'b1;
      zz_rom_62[74] = 1'b1;
      zz_rom_62[75] = 1'b1;
      zz_rom_62[76] = 1'b1;
      zz_rom_62[77] = 1'b1;
      zz_rom_62[78] = 1'b1;
      zz_rom_62[79] = 1'b1;
      zz_rom_62[80] = 1'b1;
      zz_rom_62[81] = 1'b1;
      zz_rom_62[82] = 1'b1;
      zz_rom_62[83] = 1'b1;
      zz_rom_62[84] = 1'b1;
      zz_rom_62[85] = 1'b1;
      zz_rom_62[86] = 1'b1;
      zz_rom_62[87] = 1'b1;
      zz_rom_62[88] = 1'b1;
      zz_rom_62[89] = 1'b1;
      zz_rom_62[90] = 1'b1;
      zz_rom_62[91] = 1'b1;
      zz_rom_62[92] = 1'b1;
      zz_rom_62[93] = 1'b1;
      zz_rom_62[94] = 1'b1;
      zz_rom_62[95] = 1'b1;
      zz_rom_62[96] = 1'b1;
      zz_rom_62[97] = 1'b1;
      zz_rom_62[98] = 1'b1;
      zz_rom_62[99] = 1'b0;
    end
  endfunction
  wire [99:0] _zz_63;
  function [99:0] zz_rom_63(input dummy);
    begin
      zz_rom_63[0] = 1'b0;
      zz_rom_63[1] = 1'b0;
      zz_rom_63[2] = 1'b1;
      zz_rom_63[3] = 1'b1;
      zz_rom_63[4] = 1'b1;
      zz_rom_63[5] = 1'b1;
      zz_rom_63[6] = 1'b1;
      zz_rom_63[7] = 1'b1;
      zz_rom_63[8] = 1'b1;
      zz_rom_63[9] = 1'b1;
      zz_rom_63[10] = 1'b1;
      zz_rom_63[11] = 1'b1;
      zz_rom_63[12] = 1'b1;
      zz_rom_63[13] = 1'b1;
      zz_rom_63[14] = 1'b1;
      zz_rom_63[15] = 1'b1;
      zz_rom_63[16] = 1'b1;
      zz_rom_63[17] = 1'b1;
      zz_rom_63[18] = 1'b1;
      zz_rom_63[19] = 1'b1;
      zz_rom_63[20] = 1'b1;
      zz_rom_63[21] = 1'b1;
      zz_rom_63[22] = 1'b1;
      zz_rom_63[23] = 1'b1;
      zz_rom_63[24] = 1'b1;
      zz_rom_63[25] = 1'b1;
      zz_rom_63[26] = 1'b1;
      zz_rom_63[27] = 1'b1;
      zz_rom_63[28] = 1'b1;
      zz_rom_63[29] = 1'b1;
      zz_rom_63[30] = 1'b1;
      zz_rom_63[31] = 1'b1;
      zz_rom_63[32] = 1'b1;
      zz_rom_63[33] = 1'b1;
      zz_rom_63[34] = 1'b1;
      zz_rom_63[35] = 1'b1;
      zz_rom_63[36] = 1'b1;
      zz_rom_63[37] = 1'b1;
      zz_rom_63[38] = 1'b1;
      zz_rom_63[39] = 1'b1;
      zz_rom_63[40] = 1'b1;
      zz_rom_63[41] = 1'b1;
      zz_rom_63[42] = 1'b1;
      zz_rom_63[43] = 1'b1;
      zz_rom_63[44] = 1'b1;
      zz_rom_63[45] = 1'b1;
      zz_rom_63[46] = 1'b1;
      zz_rom_63[47] = 1'b1;
      zz_rom_63[48] = 1'b1;
      zz_rom_63[49] = 1'b1;
      zz_rom_63[50] = 1'b1;
      zz_rom_63[51] = 1'b1;
      zz_rom_63[52] = 1'b1;
      zz_rom_63[53] = 1'b1;
      zz_rom_63[54] = 1'b1;
      zz_rom_63[55] = 1'b1;
      zz_rom_63[56] = 1'b1;
      zz_rom_63[57] = 1'b1;
      zz_rom_63[58] = 1'b1;
      zz_rom_63[59] = 1'b1;
      zz_rom_63[60] = 1'b1;
      zz_rom_63[61] = 1'b1;
      zz_rom_63[62] = 1'b1;
      zz_rom_63[63] = 1'b1;
      zz_rom_63[64] = 1'b1;
      zz_rom_63[65] = 1'b1;
      zz_rom_63[66] = 1'b1;
      zz_rom_63[67] = 1'b1;
      zz_rom_63[68] = 1'b1;
      zz_rom_63[69] = 1'b1;
      zz_rom_63[70] = 1'b1;
      zz_rom_63[71] = 1'b1;
      zz_rom_63[72] = 1'b1;
      zz_rom_63[73] = 1'b1;
      zz_rom_63[74] = 1'b1;
      zz_rom_63[75] = 1'b1;
      zz_rom_63[76] = 1'b1;
      zz_rom_63[77] = 1'b1;
      zz_rom_63[78] = 1'b1;
      zz_rom_63[79] = 1'b1;
      zz_rom_63[80] = 1'b1;
      zz_rom_63[81] = 1'b1;
      zz_rom_63[82] = 1'b1;
      zz_rom_63[83] = 1'b1;
      zz_rom_63[84] = 1'b1;
      zz_rom_63[85] = 1'b1;
      zz_rom_63[86] = 1'b1;
      zz_rom_63[87] = 1'b1;
      zz_rom_63[88] = 1'b1;
      zz_rom_63[89] = 1'b1;
      zz_rom_63[90] = 1'b1;
      zz_rom_63[91] = 1'b1;
      zz_rom_63[92] = 1'b1;
      zz_rom_63[93] = 1'b1;
      zz_rom_63[94] = 1'b1;
      zz_rom_63[95] = 1'b1;
      zz_rom_63[96] = 1'b1;
      zz_rom_63[97] = 1'b1;
      zz_rom_63[98] = 1'b1;
      zz_rom_63[99] = 1'b0;
    end
  endfunction
  wire [99:0] _zz_64;
  function [99:0] zz_rom_64(input dummy);
    begin
      zz_rom_64[0] = 1'b0;
      zz_rom_64[1] = 1'b0;
      zz_rom_64[2] = 1'b1;
      zz_rom_64[3] = 1'b1;
      zz_rom_64[4] = 1'b1;
      zz_rom_64[5] = 1'b1;
      zz_rom_64[6] = 1'b1;
      zz_rom_64[7] = 1'b1;
      zz_rom_64[8] = 1'b1;
      zz_rom_64[9] = 1'b1;
      zz_rom_64[10] = 1'b1;
      zz_rom_64[11] = 1'b1;
      zz_rom_64[12] = 1'b1;
      zz_rom_64[13] = 1'b1;
      zz_rom_64[14] = 1'b1;
      zz_rom_64[15] = 1'b1;
      zz_rom_64[16] = 1'b1;
      zz_rom_64[17] = 1'b1;
      zz_rom_64[18] = 1'b1;
      zz_rom_64[19] = 1'b1;
      zz_rom_64[20] = 1'b1;
      zz_rom_64[21] = 1'b1;
      zz_rom_64[22] = 1'b1;
      zz_rom_64[23] = 1'b1;
      zz_rom_64[24] = 1'b1;
      zz_rom_64[25] = 1'b1;
      zz_rom_64[26] = 1'b1;
      zz_rom_64[27] = 1'b1;
      zz_rom_64[28] = 1'b1;
      zz_rom_64[29] = 1'b1;
      zz_rom_64[30] = 1'b1;
      zz_rom_64[31] = 1'b1;
      zz_rom_64[32] = 1'b1;
      zz_rom_64[33] = 1'b1;
      zz_rom_64[34] = 1'b1;
      zz_rom_64[35] = 1'b1;
      zz_rom_64[36] = 1'b1;
      zz_rom_64[37] = 1'b1;
      zz_rom_64[38] = 1'b1;
      zz_rom_64[39] = 1'b1;
      zz_rom_64[40] = 1'b1;
      zz_rom_64[41] = 1'b1;
      zz_rom_64[42] = 1'b1;
      zz_rom_64[43] = 1'b1;
      zz_rom_64[44] = 1'b1;
      zz_rom_64[45] = 1'b1;
      zz_rom_64[46] = 1'b1;
      zz_rom_64[47] = 1'b1;
      zz_rom_64[48] = 1'b1;
      zz_rom_64[49] = 1'b1;
      zz_rom_64[50] = 1'b1;
      zz_rom_64[51] = 1'b1;
      zz_rom_64[52] = 1'b1;
      zz_rom_64[53] = 1'b1;
      zz_rom_64[54] = 1'b1;
      zz_rom_64[55] = 1'b1;
      zz_rom_64[56] = 1'b1;
      zz_rom_64[57] = 1'b1;
      zz_rom_64[58] = 1'b1;
      zz_rom_64[59] = 1'b1;
      zz_rom_64[60] = 1'b1;
      zz_rom_64[61] = 1'b1;
      zz_rom_64[62] = 1'b1;
      zz_rom_64[63] = 1'b1;
      zz_rom_64[64] = 1'b1;
      zz_rom_64[65] = 1'b1;
      zz_rom_64[66] = 1'b1;
      zz_rom_64[67] = 1'b1;
      zz_rom_64[68] = 1'b1;
      zz_rom_64[69] = 1'b1;
      zz_rom_64[70] = 1'b1;
      zz_rom_64[71] = 1'b1;
      zz_rom_64[72] = 1'b1;
      zz_rom_64[73] = 1'b1;
      zz_rom_64[74] = 1'b1;
      zz_rom_64[75] = 1'b1;
      zz_rom_64[76] = 1'b1;
      zz_rom_64[77] = 1'b1;
      zz_rom_64[78] = 1'b1;
      zz_rom_64[79] = 1'b1;
      zz_rom_64[80] = 1'b1;
      zz_rom_64[81] = 1'b1;
      zz_rom_64[82] = 1'b1;
      zz_rom_64[83] = 1'b1;
      zz_rom_64[84] = 1'b1;
      zz_rom_64[85] = 1'b1;
      zz_rom_64[86] = 1'b1;
      zz_rom_64[87] = 1'b1;
      zz_rom_64[88] = 1'b1;
      zz_rom_64[89] = 1'b1;
      zz_rom_64[90] = 1'b1;
      zz_rom_64[91] = 1'b1;
      zz_rom_64[92] = 1'b1;
      zz_rom_64[93] = 1'b1;
      zz_rom_64[94] = 1'b1;
      zz_rom_64[95] = 1'b1;
      zz_rom_64[96] = 1'b1;
      zz_rom_64[97] = 1'b1;
      zz_rom_64[98] = 1'b1;
      zz_rom_64[99] = 1'b0;
    end
  endfunction
  wire [99:0] _zz_65;
  function [99:0] zz_rom_65(input dummy);
    begin
      zz_rom_65[0] = 1'b0;
      zz_rom_65[1] = 1'b0;
      zz_rom_65[2] = 1'b0;
      zz_rom_65[3] = 1'b1;
      zz_rom_65[4] = 1'b1;
      zz_rom_65[5] = 1'b1;
      zz_rom_65[6] = 1'b1;
      zz_rom_65[7] = 1'b1;
      zz_rom_65[8] = 1'b1;
      zz_rom_65[9] = 1'b1;
      zz_rom_65[10] = 1'b1;
      zz_rom_65[11] = 1'b1;
      zz_rom_65[12] = 1'b1;
      zz_rom_65[13] = 1'b1;
      zz_rom_65[14] = 1'b1;
      zz_rom_65[15] = 1'b1;
      zz_rom_65[16] = 1'b1;
      zz_rom_65[17] = 1'b1;
      zz_rom_65[18] = 1'b1;
      zz_rom_65[19] = 1'b1;
      zz_rom_65[20] = 1'b1;
      zz_rom_65[21] = 1'b1;
      zz_rom_65[22] = 1'b1;
      zz_rom_65[23] = 1'b1;
      zz_rom_65[24] = 1'b1;
      zz_rom_65[25] = 1'b1;
      zz_rom_65[26] = 1'b1;
      zz_rom_65[27] = 1'b1;
      zz_rom_65[28] = 1'b1;
      zz_rom_65[29] = 1'b1;
      zz_rom_65[30] = 1'b1;
      zz_rom_65[31] = 1'b1;
      zz_rom_65[32] = 1'b1;
      zz_rom_65[33] = 1'b1;
      zz_rom_65[34] = 1'b1;
      zz_rom_65[35] = 1'b1;
      zz_rom_65[36] = 1'b1;
      zz_rom_65[37] = 1'b1;
      zz_rom_65[38] = 1'b1;
      zz_rom_65[39] = 1'b1;
      zz_rom_65[40] = 1'b1;
      zz_rom_65[41] = 1'b1;
      zz_rom_65[42] = 1'b1;
      zz_rom_65[43] = 1'b1;
      zz_rom_65[44] = 1'b1;
      zz_rom_65[45] = 1'b1;
      zz_rom_65[46] = 1'b1;
      zz_rom_65[47] = 1'b1;
      zz_rom_65[48] = 1'b1;
      zz_rom_65[49] = 1'b1;
      zz_rom_65[50] = 1'b1;
      zz_rom_65[51] = 1'b1;
      zz_rom_65[52] = 1'b1;
      zz_rom_65[53] = 1'b1;
      zz_rom_65[54] = 1'b1;
      zz_rom_65[55] = 1'b1;
      zz_rom_65[56] = 1'b1;
      zz_rom_65[57] = 1'b1;
      zz_rom_65[58] = 1'b1;
      zz_rom_65[59] = 1'b1;
      zz_rom_65[60] = 1'b1;
      zz_rom_65[61] = 1'b1;
      zz_rom_65[62] = 1'b1;
      zz_rom_65[63] = 1'b1;
      zz_rom_65[64] = 1'b1;
      zz_rom_65[65] = 1'b1;
      zz_rom_65[66] = 1'b1;
      zz_rom_65[67] = 1'b1;
      zz_rom_65[68] = 1'b1;
      zz_rom_65[69] = 1'b1;
      zz_rom_65[70] = 1'b1;
      zz_rom_65[71] = 1'b1;
      zz_rom_65[72] = 1'b1;
      zz_rom_65[73] = 1'b1;
      zz_rom_65[74] = 1'b1;
      zz_rom_65[75] = 1'b1;
      zz_rom_65[76] = 1'b1;
      zz_rom_65[77] = 1'b1;
      zz_rom_65[78] = 1'b1;
      zz_rom_65[79] = 1'b1;
      zz_rom_65[80] = 1'b1;
      zz_rom_65[81] = 1'b1;
      zz_rom_65[82] = 1'b1;
      zz_rom_65[83] = 1'b1;
      zz_rom_65[84] = 1'b1;
      zz_rom_65[85] = 1'b1;
      zz_rom_65[86] = 1'b1;
      zz_rom_65[87] = 1'b1;
      zz_rom_65[88] = 1'b1;
      zz_rom_65[89] = 1'b1;
      zz_rom_65[90] = 1'b1;
      zz_rom_65[91] = 1'b1;
      zz_rom_65[92] = 1'b1;
      zz_rom_65[93] = 1'b1;
      zz_rom_65[94] = 1'b1;
      zz_rom_65[95] = 1'b1;
      zz_rom_65[96] = 1'b1;
      zz_rom_65[97] = 1'b1;
      zz_rom_65[98] = 1'b0;
      zz_rom_65[99] = 1'b0;
    end
  endfunction
  wire [99:0] _zz_66;
  function [99:0] zz_rom_66(input dummy);
    begin
      zz_rom_66[0] = 1'b0;
      zz_rom_66[1] = 1'b0;
      zz_rom_66[2] = 1'b0;
      zz_rom_66[3] = 1'b1;
      zz_rom_66[4] = 1'b1;
      zz_rom_66[5] = 1'b1;
      zz_rom_66[6] = 1'b1;
      zz_rom_66[7] = 1'b1;
      zz_rom_66[8] = 1'b1;
      zz_rom_66[9] = 1'b1;
      zz_rom_66[10] = 1'b1;
      zz_rom_66[11] = 1'b1;
      zz_rom_66[12] = 1'b1;
      zz_rom_66[13] = 1'b1;
      zz_rom_66[14] = 1'b1;
      zz_rom_66[15] = 1'b1;
      zz_rom_66[16] = 1'b1;
      zz_rom_66[17] = 1'b1;
      zz_rom_66[18] = 1'b1;
      zz_rom_66[19] = 1'b1;
      zz_rom_66[20] = 1'b1;
      zz_rom_66[21] = 1'b1;
      zz_rom_66[22] = 1'b1;
      zz_rom_66[23] = 1'b1;
      zz_rom_66[24] = 1'b1;
      zz_rom_66[25] = 1'b1;
      zz_rom_66[26] = 1'b1;
      zz_rom_66[27] = 1'b1;
      zz_rom_66[28] = 1'b1;
      zz_rom_66[29] = 1'b1;
      zz_rom_66[30] = 1'b1;
      zz_rom_66[31] = 1'b1;
      zz_rom_66[32] = 1'b1;
      zz_rom_66[33] = 1'b1;
      zz_rom_66[34] = 1'b1;
      zz_rom_66[35] = 1'b1;
      zz_rom_66[36] = 1'b1;
      zz_rom_66[37] = 1'b1;
      zz_rom_66[38] = 1'b1;
      zz_rom_66[39] = 1'b1;
      zz_rom_66[40] = 1'b1;
      zz_rom_66[41] = 1'b1;
      zz_rom_66[42] = 1'b1;
      zz_rom_66[43] = 1'b1;
      zz_rom_66[44] = 1'b1;
      zz_rom_66[45] = 1'b1;
      zz_rom_66[46] = 1'b1;
      zz_rom_66[47] = 1'b1;
      zz_rom_66[48] = 1'b1;
      zz_rom_66[49] = 1'b1;
      zz_rom_66[50] = 1'b1;
      zz_rom_66[51] = 1'b1;
      zz_rom_66[52] = 1'b1;
      zz_rom_66[53] = 1'b1;
      zz_rom_66[54] = 1'b1;
      zz_rom_66[55] = 1'b1;
      zz_rom_66[56] = 1'b1;
      zz_rom_66[57] = 1'b1;
      zz_rom_66[58] = 1'b1;
      zz_rom_66[59] = 1'b1;
      zz_rom_66[60] = 1'b1;
      zz_rom_66[61] = 1'b1;
      zz_rom_66[62] = 1'b1;
      zz_rom_66[63] = 1'b1;
      zz_rom_66[64] = 1'b1;
      zz_rom_66[65] = 1'b1;
      zz_rom_66[66] = 1'b1;
      zz_rom_66[67] = 1'b1;
      zz_rom_66[68] = 1'b1;
      zz_rom_66[69] = 1'b1;
      zz_rom_66[70] = 1'b1;
      zz_rom_66[71] = 1'b1;
      zz_rom_66[72] = 1'b1;
      zz_rom_66[73] = 1'b1;
      zz_rom_66[74] = 1'b1;
      zz_rom_66[75] = 1'b1;
      zz_rom_66[76] = 1'b1;
      zz_rom_66[77] = 1'b1;
      zz_rom_66[78] = 1'b1;
      zz_rom_66[79] = 1'b1;
      zz_rom_66[80] = 1'b1;
      zz_rom_66[81] = 1'b1;
      zz_rom_66[82] = 1'b1;
      zz_rom_66[83] = 1'b1;
      zz_rom_66[84] = 1'b1;
      zz_rom_66[85] = 1'b1;
      zz_rom_66[86] = 1'b1;
      zz_rom_66[87] = 1'b1;
      zz_rom_66[88] = 1'b1;
      zz_rom_66[89] = 1'b1;
      zz_rom_66[90] = 1'b1;
      zz_rom_66[91] = 1'b1;
      zz_rom_66[92] = 1'b1;
      zz_rom_66[93] = 1'b1;
      zz_rom_66[94] = 1'b1;
      zz_rom_66[95] = 1'b1;
      zz_rom_66[96] = 1'b1;
      zz_rom_66[97] = 1'b1;
      zz_rom_66[98] = 1'b0;
      zz_rom_66[99] = 1'b0;
    end
  endfunction
  wire [99:0] _zz_67;
  function [99:0] zz_rom_67(input dummy);
    begin
      zz_rom_67[0] = 1'b0;
      zz_rom_67[1] = 1'b0;
      zz_rom_67[2] = 1'b0;
      zz_rom_67[3] = 1'b1;
      zz_rom_67[4] = 1'b1;
      zz_rom_67[5] = 1'b1;
      zz_rom_67[6] = 1'b1;
      zz_rom_67[7] = 1'b1;
      zz_rom_67[8] = 1'b1;
      zz_rom_67[9] = 1'b1;
      zz_rom_67[10] = 1'b1;
      zz_rom_67[11] = 1'b1;
      zz_rom_67[12] = 1'b1;
      zz_rom_67[13] = 1'b1;
      zz_rom_67[14] = 1'b1;
      zz_rom_67[15] = 1'b1;
      zz_rom_67[16] = 1'b1;
      zz_rom_67[17] = 1'b1;
      zz_rom_67[18] = 1'b1;
      zz_rom_67[19] = 1'b1;
      zz_rom_67[20] = 1'b1;
      zz_rom_67[21] = 1'b1;
      zz_rom_67[22] = 1'b1;
      zz_rom_67[23] = 1'b1;
      zz_rom_67[24] = 1'b1;
      zz_rom_67[25] = 1'b1;
      zz_rom_67[26] = 1'b1;
      zz_rom_67[27] = 1'b1;
      zz_rom_67[28] = 1'b1;
      zz_rom_67[29] = 1'b1;
      zz_rom_67[30] = 1'b1;
      zz_rom_67[31] = 1'b1;
      zz_rom_67[32] = 1'b1;
      zz_rom_67[33] = 1'b1;
      zz_rom_67[34] = 1'b1;
      zz_rom_67[35] = 1'b1;
      zz_rom_67[36] = 1'b1;
      zz_rom_67[37] = 1'b1;
      zz_rom_67[38] = 1'b1;
      zz_rom_67[39] = 1'b1;
      zz_rom_67[40] = 1'b1;
      zz_rom_67[41] = 1'b1;
      zz_rom_67[42] = 1'b1;
      zz_rom_67[43] = 1'b1;
      zz_rom_67[44] = 1'b1;
      zz_rom_67[45] = 1'b1;
      zz_rom_67[46] = 1'b1;
      zz_rom_67[47] = 1'b1;
      zz_rom_67[48] = 1'b1;
      zz_rom_67[49] = 1'b1;
      zz_rom_67[50] = 1'b1;
      zz_rom_67[51] = 1'b1;
      zz_rom_67[52] = 1'b1;
      zz_rom_67[53] = 1'b1;
      zz_rom_67[54] = 1'b1;
      zz_rom_67[55] = 1'b1;
      zz_rom_67[56] = 1'b1;
      zz_rom_67[57] = 1'b1;
      zz_rom_67[58] = 1'b1;
      zz_rom_67[59] = 1'b1;
      zz_rom_67[60] = 1'b1;
      zz_rom_67[61] = 1'b1;
      zz_rom_67[62] = 1'b1;
      zz_rom_67[63] = 1'b1;
      zz_rom_67[64] = 1'b1;
      zz_rom_67[65] = 1'b1;
      zz_rom_67[66] = 1'b1;
      zz_rom_67[67] = 1'b1;
      zz_rom_67[68] = 1'b1;
      zz_rom_67[69] = 1'b1;
      zz_rom_67[70] = 1'b1;
      zz_rom_67[71] = 1'b1;
      zz_rom_67[72] = 1'b1;
      zz_rom_67[73] = 1'b1;
      zz_rom_67[74] = 1'b1;
      zz_rom_67[75] = 1'b1;
      zz_rom_67[76] = 1'b1;
      zz_rom_67[77] = 1'b1;
      zz_rom_67[78] = 1'b1;
      zz_rom_67[79] = 1'b1;
      zz_rom_67[80] = 1'b1;
      zz_rom_67[81] = 1'b1;
      zz_rom_67[82] = 1'b1;
      zz_rom_67[83] = 1'b1;
      zz_rom_67[84] = 1'b1;
      zz_rom_67[85] = 1'b1;
      zz_rom_67[86] = 1'b1;
      zz_rom_67[87] = 1'b1;
      zz_rom_67[88] = 1'b1;
      zz_rom_67[89] = 1'b1;
      zz_rom_67[90] = 1'b1;
      zz_rom_67[91] = 1'b1;
      zz_rom_67[92] = 1'b1;
      zz_rom_67[93] = 1'b1;
      zz_rom_67[94] = 1'b1;
      zz_rom_67[95] = 1'b1;
      zz_rom_67[96] = 1'b1;
      zz_rom_67[97] = 1'b1;
      zz_rom_67[98] = 1'b0;
      zz_rom_67[99] = 1'b0;
    end
  endfunction
  wire [99:0] _zz_68;
  function [99:0] zz_rom_68(input dummy);
    begin
      zz_rom_68[0] = 1'b0;
      zz_rom_68[1] = 1'b0;
      zz_rom_68[2] = 1'b0;
      zz_rom_68[3] = 1'b0;
      zz_rom_68[4] = 1'b1;
      zz_rom_68[5] = 1'b1;
      zz_rom_68[6] = 1'b1;
      zz_rom_68[7] = 1'b1;
      zz_rom_68[8] = 1'b1;
      zz_rom_68[9] = 1'b1;
      zz_rom_68[10] = 1'b1;
      zz_rom_68[11] = 1'b1;
      zz_rom_68[12] = 1'b1;
      zz_rom_68[13] = 1'b1;
      zz_rom_68[14] = 1'b1;
      zz_rom_68[15] = 1'b1;
      zz_rom_68[16] = 1'b1;
      zz_rom_68[17] = 1'b1;
      zz_rom_68[18] = 1'b1;
      zz_rom_68[19] = 1'b1;
      zz_rom_68[20] = 1'b1;
      zz_rom_68[21] = 1'b1;
      zz_rom_68[22] = 1'b1;
      zz_rom_68[23] = 1'b1;
      zz_rom_68[24] = 1'b1;
      zz_rom_68[25] = 1'b1;
      zz_rom_68[26] = 1'b1;
      zz_rom_68[27] = 1'b1;
      zz_rom_68[28] = 1'b1;
      zz_rom_68[29] = 1'b1;
      zz_rom_68[30] = 1'b1;
      zz_rom_68[31] = 1'b1;
      zz_rom_68[32] = 1'b1;
      zz_rom_68[33] = 1'b1;
      zz_rom_68[34] = 1'b1;
      zz_rom_68[35] = 1'b1;
      zz_rom_68[36] = 1'b1;
      zz_rom_68[37] = 1'b1;
      zz_rom_68[38] = 1'b1;
      zz_rom_68[39] = 1'b1;
      zz_rom_68[40] = 1'b1;
      zz_rom_68[41] = 1'b1;
      zz_rom_68[42] = 1'b1;
      zz_rom_68[43] = 1'b1;
      zz_rom_68[44] = 1'b1;
      zz_rom_68[45] = 1'b1;
      zz_rom_68[46] = 1'b1;
      zz_rom_68[47] = 1'b1;
      zz_rom_68[48] = 1'b1;
      zz_rom_68[49] = 1'b1;
      zz_rom_68[50] = 1'b1;
      zz_rom_68[51] = 1'b1;
      zz_rom_68[52] = 1'b1;
      zz_rom_68[53] = 1'b1;
      zz_rom_68[54] = 1'b1;
      zz_rom_68[55] = 1'b1;
      zz_rom_68[56] = 1'b1;
      zz_rom_68[57] = 1'b1;
      zz_rom_68[58] = 1'b1;
      zz_rom_68[59] = 1'b1;
      zz_rom_68[60] = 1'b1;
      zz_rom_68[61] = 1'b1;
      zz_rom_68[62] = 1'b1;
      zz_rom_68[63] = 1'b1;
      zz_rom_68[64] = 1'b1;
      zz_rom_68[65] = 1'b1;
      zz_rom_68[66] = 1'b1;
      zz_rom_68[67] = 1'b1;
      zz_rom_68[68] = 1'b1;
      zz_rom_68[69] = 1'b1;
      zz_rom_68[70] = 1'b1;
      zz_rom_68[71] = 1'b1;
      zz_rom_68[72] = 1'b1;
      zz_rom_68[73] = 1'b1;
      zz_rom_68[74] = 1'b1;
      zz_rom_68[75] = 1'b1;
      zz_rom_68[76] = 1'b1;
      zz_rom_68[77] = 1'b1;
      zz_rom_68[78] = 1'b1;
      zz_rom_68[79] = 1'b1;
      zz_rom_68[80] = 1'b1;
      zz_rom_68[81] = 1'b1;
      zz_rom_68[82] = 1'b1;
      zz_rom_68[83] = 1'b1;
      zz_rom_68[84] = 1'b1;
      zz_rom_68[85] = 1'b1;
      zz_rom_68[86] = 1'b1;
      zz_rom_68[87] = 1'b1;
      zz_rom_68[88] = 1'b1;
      zz_rom_68[89] = 1'b1;
      zz_rom_68[90] = 1'b1;
      zz_rom_68[91] = 1'b1;
      zz_rom_68[92] = 1'b1;
      zz_rom_68[93] = 1'b1;
      zz_rom_68[94] = 1'b1;
      zz_rom_68[95] = 1'b1;
      zz_rom_68[96] = 1'b1;
      zz_rom_68[97] = 1'b0;
      zz_rom_68[98] = 1'b0;
      zz_rom_68[99] = 1'b0;
    end
  endfunction
  wire [99:0] _zz_69;
  function [99:0] zz_rom_69(input dummy);
    begin
      zz_rom_69[0] = 1'b0;
      zz_rom_69[1] = 1'b0;
      zz_rom_69[2] = 1'b0;
      zz_rom_69[3] = 1'b0;
      zz_rom_69[4] = 1'b1;
      zz_rom_69[5] = 1'b1;
      zz_rom_69[6] = 1'b1;
      zz_rom_69[7] = 1'b1;
      zz_rom_69[8] = 1'b1;
      zz_rom_69[9] = 1'b1;
      zz_rom_69[10] = 1'b1;
      zz_rom_69[11] = 1'b1;
      zz_rom_69[12] = 1'b1;
      zz_rom_69[13] = 1'b1;
      zz_rom_69[14] = 1'b1;
      zz_rom_69[15] = 1'b1;
      zz_rom_69[16] = 1'b1;
      zz_rom_69[17] = 1'b1;
      zz_rom_69[18] = 1'b1;
      zz_rom_69[19] = 1'b1;
      zz_rom_69[20] = 1'b1;
      zz_rom_69[21] = 1'b1;
      zz_rom_69[22] = 1'b1;
      zz_rom_69[23] = 1'b1;
      zz_rom_69[24] = 1'b1;
      zz_rom_69[25] = 1'b1;
      zz_rom_69[26] = 1'b1;
      zz_rom_69[27] = 1'b1;
      zz_rom_69[28] = 1'b1;
      zz_rom_69[29] = 1'b1;
      zz_rom_69[30] = 1'b1;
      zz_rom_69[31] = 1'b1;
      zz_rom_69[32] = 1'b1;
      zz_rom_69[33] = 1'b1;
      zz_rom_69[34] = 1'b1;
      zz_rom_69[35] = 1'b1;
      zz_rom_69[36] = 1'b1;
      zz_rom_69[37] = 1'b1;
      zz_rom_69[38] = 1'b1;
      zz_rom_69[39] = 1'b1;
      zz_rom_69[40] = 1'b1;
      zz_rom_69[41] = 1'b1;
      zz_rom_69[42] = 1'b1;
      zz_rom_69[43] = 1'b1;
      zz_rom_69[44] = 1'b1;
      zz_rom_69[45] = 1'b1;
      zz_rom_69[46] = 1'b1;
      zz_rom_69[47] = 1'b1;
      zz_rom_69[48] = 1'b1;
      zz_rom_69[49] = 1'b1;
      zz_rom_69[50] = 1'b1;
      zz_rom_69[51] = 1'b1;
      zz_rom_69[52] = 1'b1;
      zz_rom_69[53] = 1'b1;
      zz_rom_69[54] = 1'b1;
      zz_rom_69[55] = 1'b1;
      zz_rom_69[56] = 1'b1;
      zz_rom_69[57] = 1'b1;
      zz_rom_69[58] = 1'b1;
      zz_rom_69[59] = 1'b1;
      zz_rom_69[60] = 1'b1;
      zz_rom_69[61] = 1'b1;
      zz_rom_69[62] = 1'b1;
      zz_rom_69[63] = 1'b1;
      zz_rom_69[64] = 1'b1;
      zz_rom_69[65] = 1'b1;
      zz_rom_69[66] = 1'b1;
      zz_rom_69[67] = 1'b1;
      zz_rom_69[68] = 1'b1;
      zz_rom_69[69] = 1'b1;
      zz_rom_69[70] = 1'b1;
      zz_rom_69[71] = 1'b1;
      zz_rom_69[72] = 1'b1;
      zz_rom_69[73] = 1'b1;
      zz_rom_69[74] = 1'b1;
      zz_rom_69[75] = 1'b1;
      zz_rom_69[76] = 1'b1;
      zz_rom_69[77] = 1'b1;
      zz_rom_69[78] = 1'b1;
      zz_rom_69[79] = 1'b1;
      zz_rom_69[80] = 1'b1;
      zz_rom_69[81] = 1'b1;
      zz_rom_69[82] = 1'b1;
      zz_rom_69[83] = 1'b1;
      zz_rom_69[84] = 1'b1;
      zz_rom_69[85] = 1'b1;
      zz_rom_69[86] = 1'b1;
      zz_rom_69[87] = 1'b1;
      zz_rom_69[88] = 1'b1;
      zz_rom_69[89] = 1'b1;
      zz_rom_69[90] = 1'b1;
      zz_rom_69[91] = 1'b1;
      zz_rom_69[92] = 1'b1;
      zz_rom_69[93] = 1'b1;
      zz_rom_69[94] = 1'b1;
      zz_rom_69[95] = 1'b1;
      zz_rom_69[96] = 1'b1;
      zz_rom_69[97] = 1'b0;
      zz_rom_69[98] = 1'b0;
      zz_rom_69[99] = 1'b0;
    end
  endfunction
  wire [99:0] _zz_70;
  function [99:0] zz_rom_70(input dummy);
    begin
      zz_rom_70[0] = 1'b0;
      zz_rom_70[1] = 1'b0;
      zz_rom_70[2] = 1'b0;
      zz_rom_70[3] = 1'b0;
      zz_rom_70[4] = 1'b0;
      zz_rom_70[5] = 1'b1;
      zz_rom_70[6] = 1'b1;
      zz_rom_70[7] = 1'b1;
      zz_rom_70[8] = 1'b1;
      zz_rom_70[9] = 1'b1;
      zz_rom_70[10] = 1'b1;
      zz_rom_70[11] = 1'b1;
      zz_rom_70[12] = 1'b1;
      zz_rom_70[13] = 1'b1;
      zz_rom_70[14] = 1'b1;
      zz_rom_70[15] = 1'b1;
      zz_rom_70[16] = 1'b1;
      zz_rom_70[17] = 1'b1;
      zz_rom_70[18] = 1'b1;
      zz_rom_70[19] = 1'b1;
      zz_rom_70[20] = 1'b1;
      zz_rom_70[21] = 1'b1;
      zz_rom_70[22] = 1'b1;
      zz_rom_70[23] = 1'b1;
      zz_rom_70[24] = 1'b1;
      zz_rom_70[25] = 1'b1;
      zz_rom_70[26] = 1'b1;
      zz_rom_70[27] = 1'b1;
      zz_rom_70[28] = 1'b1;
      zz_rom_70[29] = 1'b1;
      zz_rom_70[30] = 1'b1;
      zz_rom_70[31] = 1'b1;
      zz_rom_70[32] = 1'b1;
      zz_rom_70[33] = 1'b1;
      zz_rom_70[34] = 1'b1;
      zz_rom_70[35] = 1'b1;
      zz_rom_70[36] = 1'b1;
      zz_rom_70[37] = 1'b1;
      zz_rom_70[38] = 1'b1;
      zz_rom_70[39] = 1'b1;
      zz_rom_70[40] = 1'b1;
      zz_rom_70[41] = 1'b1;
      zz_rom_70[42] = 1'b1;
      zz_rom_70[43] = 1'b1;
      zz_rom_70[44] = 1'b1;
      zz_rom_70[45] = 1'b1;
      zz_rom_70[46] = 1'b1;
      zz_rom_70[47] = 1'b1;
      zz_rom_70[48] = 1'b1;
      zz_rom_70[49] = 1'b1;
      zz_rom_70[50] = 1'b1;
      zz_rom_70[51] = 1'b1;
      zz_rom_70[52] = 1'b1;
      zz_rom_70[53] = 1'b1;
      zz_rom_70[54] = 1'b1;
      zz_rom_70[55] = 1'b1;
      zz_rom_70[56] = 1'b1;
      zz_rom_70[57] = 1'b1;
      zz_rom_70[58] = 1'b1;
      zz_rom_70[59] = 1'b1;
      zz_rom_70[60] = 1'b1;
      zz_rom_70[61] = 1'b1;
      zz_rom_70[62] = 1'b1;
      zz_rom_70[63] = 1'b1;
      zz_rom_70[64] = 1'b1;
      zz_rom_70[65] = 1'b1;
      zz_rom_70[66] = 1'b1;
      zz_rom_70[67] = 1'b1;
      zz_rom_70[68] = 1'b1;
      zz_rom_70[69] = 1'b1;
      zz_rom_70[70] = 1'b1;
      zz_rom_70[71] = 1'b1;
      zz_rom_70[72] = 1'b1;
      zz_rom_70[73] = 1'b1;
      zz_rom_70[74] = 1'b1;
      zz_rom_70[75] = 1'b1;
      zz_rom_70[76] = 1'b1;
      zz_rom_70[77] = 1'b1;
      zz_rom_70[78] = 1'b1;
      zz_rom_70[79] = 1'b1;
      zz_rom_70[80] = 1'b1;
      zz_rom_70[81] = 1'b1;
      zz_rom_70[82] = 1'b1;
      zz_rom_70[83] = 1'b1;
      zz_rom_70[84] = 1'b1;
      zz_rom_70[85] = 1'b1;
      zz_rom_70[86] = 1'b1;
      zz_rom_70[87] = 1'b1;
      zz_rom_70[88] = 1'b1;
      zz_rom_70[89] = 1'b1;
      zz_rom_70[90] = 1'b1;
      zz_rom_70[91] = 1'b1;
      zz_rom_70[92] = 1'b1;
      zz_rom_70[93] = 1'b1;
      zz_rom_70[94] = 1'b1;
      zz_rom_70[95] = 1'b1;
      zz_rom_70[96] = 1'b0;
      zz_rom_70[97] = 1'b0;
      zz_rom_70[98] = 1'b0;
      zz_rom_70[99] = 1'b0;
    end
  endfunction
  wire [99:0] _zz_71;
  function [99:0] zz_rom_71(input dummy);
    begin
      zz_rom_71[0] = 1'b0;
      zz_rom_71[1] = 1'b0;
      zz_rom_71[2] = 1'b0;
      zz_rom_71[3] = 1'b0;
      zz_rom_71[4] = 1'b0;
      zz_rom_71[5] = 1'b1;
      zz_rom_71[6] = 1'b1;
      zz_rom_71[7] = 1'b1;
      zz_rom_71[8] = 1'b1;
      zz_rom_71[9] = 1'b1;
      zz_rom_71[10] = 1'b1;
      zz_rom_71[11] = 1'b1;
      zz_rom_71[12] = 1'b1;
      zz_rom_71[13] = 1'b1;
      zz_rom_71[14] = 1'b1;
      zz_rom_71[15] = 1'b1;
      zz_rom_71[16] = 1'b1;
      zz_rom_71[17] = 1'b1;
      zz_rom_71[18] = 1'b1;
      zz_rom_71[19] = 1'b1;
      zz_rom_71[20] = 1'b1;
      zz_rom_71[21] = 1'b1;
      zz_rom_71[22] = 1'b1;
      zz_rom_71[23] = 1'b1;
      zz_rom_71[24] = 1'b1;
      zz_rom_71[25] = 1'b1;
      zz_rom_71[26] = 1'b1;
      zz_rom_71[27] = 1'b1;
      zz_rom_71[28] = 1'b1;
      zz_rom_71[29] = 1'b1;
      zz_rom_71[30] = 1'b1;
      zz_rom_71[31] = 1'b1;
      zz_rom_71[32] = 1'b1;
      zz_rom_71[33] = 1'b1;
      zz_rom_71[34] = 1'b1;
      zz_rom_71[35] = 1'b1;
      zz_rom_71[36] = 1'b1;
      zz_rom_71[37] = 1'b1;
      zz_rom_71[38] = 1'b1;
      zz_rom_71[39] = 1'b1;
      zz_rom_71[40] = 1'b1;
      zz_rom_71[41] = 1'b1;
      zz_rom_71[42] = 1'b1;
      zz_rom_71[43] = 1'b1;
      zz_rom_71[44] = 1'b1;
      zz_rom_71[45] = 1'b1;
      zz_rom_71[46] = 1'b1;
      zz_rom_71[47] = 1'b1;
      zz_rom_71[48] = 1'b1;
      zz_rom_71[49] = 1'b1;
      zz_rom_71[50] = 1'b1;
      zz_rom_71[51] = 1'b1;
      zz_rom_71[52] = 1'b1;
      zz_rom_71[53] = 1'b1;
      zz_rom_71[54] = 1'b1;
      zz_rom_71[55] = 1'b1;
      zz_rom_71[56] = 1'b1;
      zz_rom_71[57] = 1'b1;
      zz_rom_71[58] = 1'b1;
      zz_rom_71[59] = 1'b1;
      zz_rom_71[60] = 1'b1;
      zz_rom_71[61] = 1'b1;
      zz_rom_71[62] = 1'b1;
      zz_rom_71[63] = 1'b1;
      zz_rom_71[64] = 1'b1;
      zz_rom_71[65] = 1'b1;
      zz_rom_71[66] = 1'b1;
      zz_rom_71[67] = 1'b1;
      zz_rom_71[68] = 1'b1;
      zz_rom_71[69] = 1'b1;
      zz_rom_71[70] = 1'b1;
      zz_rom_71[71] = 1'b1;
      zz_rom_71[72] = 1'b1;
      zz_rom_71[73] = 1'b1;
      zz_rom_71[74] = 1'b1;
      zz_rom_71[75] = 1'b1;
      zz_rom_71[76] = 1'b1;
      zz_rom_71[77] = 1'b1;
      zz_rom_71[78] = 1'b1;
      zz_rom_71[79] = 1'b1;
      zz_rom_71[80] = 1'b1;
      zz_rom_71[81] = 1'b1;
      zz_rom_71[82] = 1'b1;
      zz_rom_71[83] = 1'b1;
      zz_rom_71[84] = 1'b1;
      zz_rom_71[85] = 1'b1;
      zz_rom_71[86] = 1'b1;
      zz_rom_71[87] = 1'b1;
      zz_rom_71[88] = 1'b1;
      zz_rom_71[89] = 1'b1;
      zz_rom_71[90] = 1'b1;
      zz_rom_71[91] = 1'b1;
      zz_rom_71[92] = 1'b1;
      zz_rom_71[93] = 1'b1;
      zz_rom_71[94] = 1'b1;
      zz_rom_71[95] = 1'b1;
      zz_rom_71[96] = 1'b0;
      zz_rom_71[97] = 1'b0;
      zz_rom_71[98] = 1'b0;
      zz_rom_71[99] = 1'b0;
    end
  endfunction
  wire [99:0] _zz_72;
  function [99:0] zz_rom_72(input dummy);
    begin
      zz_rom_72[0] = 1'b0;
      zz_rom_72[1] = 1'b0;
      zz_rom_72[2] = 1'b0;
      zz_rom_72[3] = 1'b0;
      zz_rom_72[4] = 1'b0;
      zz_rom_72[5] = 1'b0;
      zz_rom_72[6] = 1'b1;
      zz_rom_72[7] = 1'b1;
      zz_rom_72[8] = 1'b1;
      zz_rom_72[9] = 1'b1;
      zz_rom_72[10] = 1'b1;
      zz_rom_72[11] = 1'b1;
      zz_rom_72[12] = 1'b1;
      zz_rom_72[13] = 1'b1;
      zz_rom_72[14] = 1'b1;
      zz_rom_72[15] = 1'b1;
      zz_rom_72[16] = 1'b1;
      zz_rom_72[17] = 1'b1;
      zz_rom_72[18] = 1'b1;
      zz_rom_72[19] = 1'b1;
      zz_rom_72[20] = 1'b1;
      zz_rom_72[21] = 1'b1;
      zz_rom_72[22] = 1'b1;
      zz_rom_72[23] = 1'b1;
      zz_rom_72[24] = 1'b1;
      zz_rom_72[25] = 1'b1;
      zz_rom_72[26] = 1'b1;
      zz_rom_72[27] = 1'b1;
      zz_rom_72[28] = 1'b1;
      zz_rom_72[29] = 1'b1;
      zz_rom_72[30] = 1'b1;
      zz_rom_72[31] = 1'b1;
      zz_rom_72[32] = 1'b1;
      zz_rom_72[33] = 1'b1;
      zz_rom_72[34] = 1'b1;
      zz_rom_72[35] = 1'b1;
      zz_rom_72[36] = 1'b1;
      zz_rom_72[37] = 1'b1;
      zz_rom_72[38] = 1'b1;
      zz_rom_72[39] = 1'b1;
      zz_rom_72[40] = 1'b1;
      zz_rom_72[41] = 1'b1;
      zz_rom_72[42] = 1'b1;
      zz_rom_72[43] = 1'b1;
      zz_rom_72[44] = 1'b1;
      zz_rom_72[45] = 1'b1;
      zz_rom_72[46] = 1'b1;
      zz_rom_72[47] = 1'b1;
      zz_rom_72[48] = 1'b1;
      zz_rom_72[49] = 1'b1;
      zz_rom_72[50] = 1'b1;
      zz_rom_72[51] = 1'b1;
      zz_rom_72[52] = 1'b1;
      zz_rom_72[53] = 1'b1;
      zz_rom_72[54] = 1'b1;
      zz_rom_72[55] = 1'b1;
      zz_rom_72[56] = 1'b1;
      zz_rom_72[57] = 1'b1;
      zz_rom_72[58] = 1'b1;
      zz_rom_72[59] = 1'b1;
      zz_rom_72[60] = 1'b1;
      zz_rom_72[61] = 1'b1;
      zz_rom_72[62] = 1'b1;
      zz_rom_72[63] = 1'b1;
      zz_rom_72[64] = 1'b1;
      zz_rom_72[65] = 1'b1;
      zz_rom_72[66] = 1'b1;
      zz_rom_72[67] = 1'b1;
      zz_rom_72[68] = 1'b1;
      zz_rom_72[69] = 1'b1;
      zz_rom_72[70] = 1'b1;
      zz_rom_72[71] = 1'b1;
      zz_rom_72[72] = 1'b1;
      zz_rom_72[73] = 1'b1;
      zz_rom_72[74] = 1'b1;
      zz_rom_72[75] = 1'b1;
      zz_rom_72[76] = 1'b1;
      zz_rom_72[77] = 1'b1;
      zz_rom_72[78] = 1'b1;
      zz_rom_72[79] = 1'b1;
      zz_rom_72[80] = 1'b1;
      zz_rom_72[81] = 1'b1;
      zz_rom_72[82] = 1'b1;
      zz_rom_72[83] = 1'b1;
      zz_rom_72[84] = 1'b1;
      zz_rom_72[85] = 1'b1;
      zz_rom_72[86] = 1'b1;
      zz_rom_72[87] = 1'b1;
      zz_rom_72[88] = 1'b1;
      zz_rom_72[89] = 1'b1;
      zz_rom_72[90] = 1'b1;
      zz_rom_72[91] = 1'b1;
      zz_rom_72[92] = 1'b1;
      zz_rom_72[93] = 1'b1;
      zz_rom_72[94] = 1'b1;
      zz_rom_72[95] = 1'b0;
      zz_rom_72[96] = 1'b0;
      zz_rom_72[97] = 1'b0;
      zz_rom_72[98] = 1'b0;
      zz_rom_72[99] = 1'b0;
    end
  endfunction
  wire [99:0] _zz_73;
  function [99:0] zz_rom_73(input dummy);
    begin
      zz_rom_73[0] = 1'b0;
      zz_rom_73[1] = 1'b0;
      zz_rom_73[2] = 1'b0;
      zz_rom_73[3] = 1'b0;
      zz_rom_73[4] = 1'b0;
      zz_rom_73[5] = 1'b0;
      zz_rom_73[6] = 1'b1;
      zz_rom_73[7] = 1'b1;
      zz_rom_73[8] = 1'b1;
      zz_rom_73[9] = 1'b1;
      zz_rom_73[10] = 1'b1;
      zz_rom_73[11] = 1'b1;
      zz_rom_73[12] = 1'b1;
      zz_rom_73[13] = 1'b1;
      zz_rom_73[14] = 1'b1;
      zz_rom_73[15] = 1'b1;
      zz_rom_73[16] = 1'b1;
      zz_rom_73[17] = 1'b1;
      zz_rom_73[18] = 1'b1;
      zz_rom_73[19] = 1'b1;
      zz_rom_73[20] = 1'b1;
      zz_rom_73[21] = 1'b1;
      zz_rom_73[22] = 1'b1;
      zz_rom_73[23] = 1'b1;
      zz_rom_73[24] = 1'b1;
      zz_rom_73[25] = 1'b1;
      zz_rom_73[26] = 1'b1;
      zz_rom_73[27] = 1'b1;
      zz_rom_73[28] = 1'b1;
      zz_rom_73[29] = 1'b1;
      zz_rom_73[30] = 1'b1;
      zz_rom_73[31] = 1'b1;
      zz_rom_73[32] = 1'b1;
      zz_rom_73[33] = 1'b1;
      zz_rom_73[34] = 1'b1;
      zz_rom_73[35] = 1'b1;
      zz_rom_73[36] = 1'b1;
      zz_rom_73[37] = 1'b1;
      zz_rom_73[38] = 1'b1;
      zz_rom_73[39] = 1'b1;
      zz_rom_73[40] = 1'b1;
      zz_rom_73[41] = 1'b1;
      zz_rom_73[42] = 1'b1;
      zz_rom_73[43] = 1'b1;
      zz_rom_73[44] = 1'b1;
      zz_rom_73[45] = 1'b1;
      zz_rom_73[46] = 1'b1;
      zz_rom_73[47] = 1'b1;
      zz_rom_73[48] = 1'b1;
      zz_rom_73[49] = 1'b1;
      zz_rom_73[50] = 1'b1;
      zz_rom_73[51] = 1'b1;
      zz_rom_73[52] = 1'b1;
      zz_rom_73[53] = 1'b1;
      zz_rom_73[54] = 1'b1;
      zz_rom_73[55] = 1'b1;
      zz_rom_73[56] = 1'b1;
      zz_rom_73[57] = 1'b1;
      zz_rom_73[58] = 1'b1;
      zz_rom_73[59] = 1'b1;
      zz_rom_73[60] = 1'b1;
      zz_rom_73[61] = 1'b1;
      zz_rom_73[62] = 1'b1;
      zz_rom_73[63] = 1'b1;
      zz_rom_73[64] = 1'b1;
      zz_rom_73[65] = 1'b1;
      zz_rom_73[66] = 1'b1;
      zz_rom_73[67] = 1'b1;
      zz_rom_73[68] = 1'b1;
      zz_rom_73[69] = 1'b1;
      zz_rom_73[70] = 1'b1;
      zz_rom_73[71] = 1'b1;
      zz_rom_73[72] = 1'b1;
      zz_rom_73[73] = 1'b1;
      zz_rom_73[74] = 1'b1;
      zz_rom_73[75] = 1'b1;
      zz_rom_73[76] = 1'b1;
      zz_rom_73[77] = 1'b1;
      zz_rom_73[78] = 1'b1;
      zz_rom_73[79] = 1'b1;
      zz_rom_73[80] = 1'b1;
      zz_rom_73[81] = 1'b1;
      zz_rom_73[82] = 1'b1;
      zz_rom_73[83] = 1'b1;
      zz_rom_73[84] = 1'b1;
      zz_rom_73[85] = 1'b1;
      zz_rom_73[86] = 1'b1;
      zz_rom_73[87] = 1'b1;
      zz_rom_73[88] = 1'b1;
      zz_rom_73[89] = 1'b1;
      zz_rom_73[90] = 1'b1;
      zz_rom_73[91] = 1'b1;
      zz_rom_73[92] = 1'b1;
      zz_rom_73[93] = 1'b1;
      zz_rom_73[94] = 1'b1;
      zz_rom_73[95] = 1'b0;
      zz_rom_73[96] = 1'b0;
      zz_rom_73[97] = 1'b0;
      zz_rom_73[98] = 1'b0;
      zz_rom_73[99] = 1'b0;
    end
  endfunction
  wire [99:0] _zz_74;
  function [99:0] zz_rom_74(input dummy);
    begin
      zz_rom_74[0] = 1'b0;
      zz_rom_74[1] = 1'b0;
      zz_rom_74[2] = 1'b0;
      zz_rom_74[3] = 1'b0;
      zz_rom_74[4] = 1'b0;
      zz_rom_74[5] = 1'b0;
      zz_rom_74[6] = 1'b0;
      zz_rom_74[7] = 1'b1;
      zz_rom_74[8] = 1'b1;
      zz_rom_74[9] = 1'b1;
      zz_rom_74[10] = 1'b1;
      zz_rom_74[11] = 1'b1;
      zz_rom_74[12] = 1'b1;
      zz_rom_74[13] = 1'b1;
      zz_rom_74[14] = 1'b1;
      zz_rom_74[15] = 1'b1;
      zz_rom_74[16] = 1'b1;
      zz_rom_74[17] = 1'b1;
      zz_rom_74[18] = 1'b1;
      zz_rom_74[19] = 1'b1;
      zz_rom_74[20] = 1'b1;
      zz_rom_74[21] = 1'b1;
      zz_rom_74[22] = 1'b1;
      zz_rom_74[23] = 1'b1;
      zz_rom_74[24] = 1'b1;
      zz_rom_74[25] = 1'b1;
      zz_rom_74[26] = 1'b1;
      zz_rom_74[27] = 1'b1;
      zz_rom_74[28] = 1'b1;
      zz_rom_74[29] = 1'b1;
      zz_rom_74[30] = 1'b1;
      zz_rom_74[31] = 1'b1;
      zz_rom_74[32] = 1'b1;
      zz_rom_74[33] = 1'b1;
      zz_rom_74[34] = 1'b1;
      zz_rom_74[35] = 1'b1;
      zz_rom_74[36] = 1'b1;
      zz_rom_74[37] = 1'b1;
      zz_rom_74[38] = 1'b1;
      zz_rom_74[39] = 1'b1;
      zz_rom_74[40] = 1'b1;
      zz_rom_74[41] = 1'b1;
      zz_rom_74[42] = 1'b1;
      zz_rom_74[43] = 1'b1;
      zz_rom_74[44] = 1'b1;
      zz_rom_74[45] = 1'b1;
      zz_rom_74[46] = 1'b1;
      zz_rom_74[47] = 1'b1;
      zz_rom_74[48] = 1'b1;
      zz_rom_74[49] = 1'b1;
      zz_rom_74[50] = 1'b1;
      zz_rom_74[51] = 1'b1;
      zz_rom_74[52] = 1'b1;
      zz_rom_74[53] = 1'b1;
      zz_rom_74[54] = 1'b1;
      zz_rom_74[55] = 1'b1;
      zz_rom_74[56] = 1'b1;
      zz_rom_74[57] = 1'b1;
      zz_rom_74[58] = 1'b1;
      zz_rom_74[59] = 1'b1;
      zz_rom_74[60] = 1'b1;
      zz_rom_74[61] = 1'b1;
      zz_rom_74[62] = 1'b1;
      zz_rom_74[63] = 1'b1;
      zz_rom_74[64] = 1'b1;
      zz_rom_74[65] = 1'b1;
      zz_rom_74[66] = 1'b1;
      zz_rom_74[67] = 1'b1;
      zz_rom_74[68] = 1'b1;
      zz_rom_74[69] = 1'b1;
      zz_rom_74[70] = 1'b1;
      zz_rom_74[71] = 1'b1;
      zz_rom_74[72] = 1'b1;
      zz_rom_74[73] = 1'b1;
      zz_rom_74[74] = 1'b1;
      zz_rom_74[75] = 1'b1;
      zz_rom_74[76] = 1'b1;
      zz_rom_74[77] = 1'b1;
      zz_rom_74[78] = 1'b1;
      zz_rom_74[79] = 1'b1;
      zz_rom_74[80] = 1'b1;
      zz_rom_74[81] = 1'b1;
      zz_rom_74[82] = 1'b1;
      zz_rom_74[83] = 1'b1;
      zz_rom_74[84] = 1'b1;
      zz_rom_74[85] = 1'b1;
      zz_rom_74[86] = 1'b1;
      zz_rom_74[87] = 1'b1;
      zz_rom_74[88] = 1'b1;
      zz_rom_74[89] = 1'b1;
      zz_rom_74[90] = 1'b1;
      zz_rom_74[91] = 1'b1;
      zz_rom_74[92] = 1'b1;
      zz_rom_74[93] = 1'b1;
      zz_rom_74[94] = 1'b0;
      zz_rom_74[95] = 1'b0;
      zz_rom_74[96] = 1'b0;
      zz_rom_74[97] = 1'b0;
      zz_rom_74[98] = 1'b0;
      zz_rom_74[99] = 1'b0;
    end
  endfunction
  wire [99:0] _zz_75;
  function [99:0] zz_rom_75(input dummy);
    begin
      zz_rom_75[0] = 1'b0;
      zz_rom_75[1] = 1'b0;
      zz_rom_75[2] = 1'b0;
      zz_rom_75[3] = 1'b0;
      zz_rom_75[4] = 1'b0;
      zz_rom_75[5] = 1'b0;
      zz_rom_75[6] = 1'b0;
      zz_rom_75[7] = 1'b1;
      zz_rom_75[8] = 1'b1;
      zz_rom_75[9] = 1'b1;
      zz_rom_75[10] = 1'b1;
      zz_rom_75[11] = 1'b1;
      zz_rom_75[12] = 1'b1;
      zz_rom_75[13] = 1'b1;
      zz_rom_75[14] = 1'b1;
      zz_rom_75[15] = 1'b1;
      zz_rom_75[16] = 1'b1;
      zz_rom_75[17] = 1'b1;
      zz_rom_75[18] = 1'b1;
      zz_rom_75[19] = 1'b1;
      zz_rom_75[20] = 1'b1;
      zz_rom_75[21] = 1'b1;
      zz_rom_75[22] = 1'b1;
      zz_rom_75[23] = 1'b1;
      zz_rom_75[24] = 1'b1;
      zz_rom_75[25] = 1'b1;
      zz_rom_75[26] = 1'b1;
      zz_rom_75[27] = 1'b1;
      zz_rom_75[28] = 1'b1;
      zz_rom_75[29] = 1'b1;
      zz_rom_75[30] = 1'b1;
      zz_rom_75[31] = 1'b1;
      zz_rom_75[32] = 1'b1;
      zz_rom_75[33] = 1'b1;
      zz_rom_75[34] = 1'b1;
      zz_rom_75[35] = 1'b1;
      zz_rom_75[36] = 1'b1;
      zz_rom_75[37] = 1'b1;
      zz_rom_75[38] = 1'b1;
      zz_rom_75[39] = 1'b1;
      zz_rom_75[40] = 1'b1;
      zz_rom_75[41] = 1'b1;
      zz_rom_75[42] = 1'b1;
      zz_rom_75[43] = 1'b1;
      zz_rom_75[44] = 1'b1;
      zz_rom_75[45] = 1'b1;
      zz_rom_75[46] = 1'b1;
      zz_rom_75[47] = 1'b1;
      zz_rom_75[48] = 1'b1;
      zz_rom_75[49] = 1'b1;
      zz_rom_75[50] = 1'b1;
      zz_rom_75[51] = 1'b1;
      zz_rom_75[52] = 1'b1;
      zz_rom_75[53] = 1'b1;
      zz_rom_75[54] = 1'b1;
      zz_rom_75[55] = 1'b1;
      zz_rom_75[56] = 1'b1;
      zz_rom_75[57] = 1'b1;
      zz_rom_75[58] = 1'b1;
      zz_rom_75[59] = 1'b1;
      zz_rom_75[60] = 1'b1;
      zz_rom_75[61] = 1'b1;
      zz_rom_75[62] = 1'b1;
      zz_rom_75[63] = 1'b1;
      zz_rom_75[64] = 1'b1;
      zz_rom_75[65] = 1'b1;
      zz_rom_75[66] = 1'b1;
      zz_rom_75[67] = 1'b1;
      zz_rom_75[68] = 1'b1;
      zz_rom_75[69] = 1'b1;
      zz_rom_75[70] = 1'b1;
      zz_rom_75[71] = 1'b1;
      zz_rom_75[72] = 1'b1;
      zz_rom_75[73] = 1'b1;
      zz_rom_75[74] = 1'b1;
      zz_rom_75[75] = 1'b1;
      zz_rom_75[76] = 1'b1;
      zz_rom_75[77] = 1'b1;
      zz_rom_75[78] = 1'b1;
      zz_rom_75[79] = 1'b1;
      zz_rom_75[80] = 1'b1;
      zz_rom_75[81] = 1'b1;
      zz_rom_75[82] = 1'b1;
      zz_rom_75[83] = 1'b1;
      zz_rom_75[84] = 1'b1;
      zz_rom_75[85] = 1'b1;
      zz_rom_75[86] = 1'b1;
      zz_rom_75[87] = 1'b1;
      zz_rom_75[88] = 1'b1;
      zz_rom_75[89] = 1'b1;
      zz_rom_75[90] = 1'b1;
      zz_rom_75[91] = 1'b1;
      zz_rom_75[92] = 1'b1;
      zz_rom_75[93] = 1'b1;
      zz_rom_75[94] = 1'b0;
      zz_rom_75[95] = 1'b0;
      zz_rom_75[96] = 1'b0;
      zz_rom_75[97] = 1'b0;
      zz_rom_75[98] = 1'b0;
      zz_rom_75[99] = 1'b0;
    end
  endfunction
  wire [99:0] _zz_76;
  function [99:0] zz_rom_76(input dummy);
    begin
      zz_rom_76[0] = 1'b0;
      zz_rom_76[1] = 1'b0;
      zz_rom_76[2] = 1'b0;
      zz_rom_76[3] = 1'b0;
      zz_rom_76[4] = 1'b0;
      zz_rom_76[5] = 1'b0;
      zz_rom_76[6] = 1'b0;
      zz_rom_76[7] = 1'b0;
      zz_rom_76[8] = 1'b1;
      zz_rom_76[9] = 1'b1;
      zz_rom_76[10] = 1'b1;
      zz_rom_76[11] = 1'b1;
      zz_rom_76[12] = 1'b1;
      zz_rom_76[13] = 1'b1;
      zz_rom_76[14] = 1'b1;
      zz_rom_76[15] = 1'b1;
      zz_rom_76[16] = 1'b1;
      zz_rom_76[17] = 1'b1;
      zz_rom_76[18] = 1'b1;
      zz_rom_76[19] = 1'b1;
      zz_rom_76[20] = 1'b1;
      zz_rom_76[21] = 1'b1;
      zz_rom_76[22] = 1'b1;
      zz_rom_76[23] = 1'b1;
      zz_rom_76[24] = 1'b1;
      zz_rom_76[25] = 1'b1;
      zz_rom_76[26] = 1'b1;
      zz_rom_76[27] = 1'b1;
      zz_rom_76[28] = 1'b1;
      zz_rom_76[29] = 1'b1;
      zz_rom_76[30] = 1'b1;
      zz_rom_76[31] = 1'b1;
      zz_rom_76[32] = 1'b1;
      zz_rom_76[33] = 1'b1;
      zz_rom_76[34] = 1'b1;
      zz_rom_76[35] = 1'b1;
      zz_rom_76[36] = 1'b1;
      zz_rom_76[37] = 1'b1;
      zz_rom_76[38] = 1'b1;
      zz_rom_76[39] = 1'b1;
      zz_rom_76[40] = 1'b1;
      zz_rom_76[41] = 1'b1;
      zz_rom_76[42] = 1'b1;
      zz_rom_76[43] = 1'b1;
      zz_rom_76[44] = 1'b1;
      zz_rom_76[45] = 1'b1;
      zz_rom_76[46] = 1'b1;
      zz_rom_76[47] = 1'b1;
      zz_rom_76[48] = 1'b1;
      zz_rom_76[49] = 1'b1;
      zz_rom_76[50] = 1'b1;
      zz_rom_76[51] = 1'b1;
      zz_rom_76[52] = 1'b1;
      zz_rom_76[53] = 1'b1;
      zz_rom_76[54] = 1'b1;
      zz_rom_76[55] = 1'b1;
      zz_rom_76[56] = 1'b1;
      zz_rom_76[57] = 1'b1;
      zz_rom_76[58] = 1'b1;
      zz_rom_76[59] = 1'b1;
      zz_rom_76[60] = 1'b1;
      zz_rom_76[61] = 1'b1;
      zz_rom_76[62] = 1'b1;
      zz_rom_76[63] = 1'b1;
      zz_rom_76[64] = 1'b1;
      zz_rom_76[65] = 1'b1;
      zz_rom_76[66] = 1'b1;
      zz_rom_76[67] = 1'b1;
      zz_rom_76[68] = 1'b1;
      zz_rom_76[69] = 1'b1;
      zz_rom_76[70] = 1'b1;
      zz_rom_76[71] = 1'b1;
      zz_rom_76[72] = 1'b1;
      zz_rom_76[73] = 1'b1;
      zz_rom_76[74] = 1'b1;
      zz_rom_76[75] = 1'b1;
      zz_rom_76[76] = 1'b1;
      zz_rom_76[77] = 1'b1;
      zz_rom_76[78] = 1'b1;
      zz_rom_76[79] = 1'b1;
      zz_rom_76[80] = 1'b1;
      zz_rom_76[81] = 1'b1;
      zz_rom_76[82] = 1'b1;
      zz_rom_76[83] = 1'b1;
      zz_rom_76[84] = 1'b1;
      zz_rom_76[85] = 1'b1;
      zz_rom_76[86] = 1'b1;
      zz_rom_76[87] = 1'b1;
      zz_rom_76[88] = 1'b1;
      zz_rom_76[89] = 1'b1;
      zz_rom_76[90] = 1'b1;
      zz_rom_76[91] = 1'b1;
      zz_rom_76[92] = 1'b1;
      zz_rom_76[93] = 1'b0;
      zz_rom_76[94] = 1'b0;
      zz_rom_76[95] = 1'b0;
      zz_rom_76[96] = 1'b0;
      zz_rom_76[97] = 1'b0;
      zz_rom_76[98] = 1'b0;
      zz_rom_76[99] = 1'b0;
    end
  endfunction
  wire [99:0] _zz_77;
  function [99:0] zz_rom_77(input dummy);
    begin
      zz_rom_77[0] = 1'b0;
      zz_rom_77[1] = 1'b0;
      zz_rom_77[2] = 1'b0;
      zz_rom_77[3] = 1'b0;
      zz_rom_77[4] = 1'b0;
      zz_rom_77[5] = 1'b0;
      zz_rom_77[6] = 1'b0;
      zz_rom_77[7] = 1'b0;
      zz_rom_77[8] = 1'b1;
      zz_rom_77[9] = 1'b1;
      zz_rom_77[10] = 1'b1;
      zz_rom_77[11] = 1'b1;
      zz_rom_77[12] = 1'b1;
      zz_rom_77[13] = 1'b1;
      zz_rom_77[14] = 1'b1;
      zz_rom_77[15] = 1'b1;
      zz_rom_77[16] = 1'b1;
      zz_rom_77[17] = 1'b1;
      zz_rom_77[18] = 1'b1;
      zz_rom_77[19] = 1'b1;
      zz_rom_77[20] = 1'b1;
      zz_rom_77[21] = 1'b1;
      zz_rom_77[22] = 1'b1;
      zz_rom_77[23] = 1'b1;
      zz_rom_77[24] = 1'b1;
      zz_rom_77[25] = 1'b1;
      zz_rom_77[26] = 1'b1;
      zz_rom_77[27] = 1'b1;
      zz_rom_77[28] = 1'b1;
      zz_rom_77[29] = 1'b1;
      zz_rom_77[30] = 1'b1;
      zz_rom_77[31] = 1'b1;
      zz_rom_77[32] = 1'b1;
      zz_rom_77[33] = 1'b1;
      zz_rom_77[34] = 1'b1;
      zz_rom_77[35] = 1'b1;
      zz_rom_77[36] = 1'b1;
      zz_rom_77[37] = 1'b1;
      zz_rom_77[38] = 1'b1;
      zz_rom_77[39] = 1'b1;
      zz_rom_77[40] = 1'b1;
      zz_rom_77[41] = 1'b1;
      zz_rom_77[42] = 1'b1;
      zz_rom_77[43] = 1'b1;
      zz_rom_77[44] = 1'b1;
      zz_rom_77[45] = 1'b1;
      zz_rom_77[46] = 1'b1;
      zz_rom_77[47] = 1'b1;
      zz_rom_77[48] = 1'b1;
      zz_rom_77[49] = 1'b1;
      zz_rom_77[50] = 1'b1;
      zz_rom_77[51] = 1'b1;
      zz_rom_77[52] = 1'b1;
      zz_rom_77[53] = 1'b1;
      zz_rom_77[54] = 1'b1;
      zz_rom_77[55] = 1'b1;
      zz_rom_77[56] = 1'b1;
      zz_rom_77[57] = 1'b1;
      zz_rom_77[58] = 1'b1;
      zz_rom_77[59] = 1'b1;
      zz_rom_77[60] = 1'b1;
      zz_rom_77[61] = 1'b1;
      zz_rom_77[62] = 1'b1;
      zz_rom_77[63] = 1'b1;
      zz_rom_77[64] = 1'b1;
      zz_rom_77[65] = 1'b1;
      zz_rom_77[66] = 1'b1;
      zz_rom_77[67] = 1'b1;
      zz_rom_77[68] = 1'b1;
      zz_rom_77[69] = 1'b1;
      zz_rom_77[70] = 1'b1;
      zz_rom_77[71] = 1'b1;
      zz_rom_77[72] = 1'b1;
      zz_rom_77[73] = 1'b1;
      zz_rom_77[74] = 1'b1;
      zz_rom_77[75] = 1'b1;
      zz_rom_77[76] = 1'b1;
      zz_rom_77[77] = 1'b1;
      zz_rom_77[78] = 1'b1;
      zz_rom_77[79] = 1'b1;
      zz_rom_77[80] = 1'b1;
      zz_rom_77[81] = 1'b1;
      zz_rom_77[82] = 1'b1;
      zz_rom_77[83] = 1'b1;
      zz_rom_77[84] = 1'b1;
      zz_rom_77[85] = 1'b1;
      zz_rom_77[86] = 1'b1;
      zz_rom_77[87] = 1'b1;
      zz_rom_77[88] = 1'b1;
      zz_rom_77[89] = 1'b1;
      zz_rom_77[90] = 1'b1;
      zz_rom_77[91] = 1'b1;
      zz_rom_77[92] = 1'b1;
      zz_rom_77[93] = 1'b0;
      zz_rom_77[94] = 1'b0;
      zz_rom_77[95] = 1'b0;
      zz_rom_77[96] = 1'b0;
      zz_rom_77[97] = 1'b0;
      zz_rom_77[98] = 1'b0;
      zz_rom_77[99] = 1'b0;
    end
  endfunction
  wire [99:0] _zz_78;
  function [99:0] zz_rom_78(input dummy);
    begin
      zz_rom_78[0] = 1'b0;
      zz_rom_78[1] = 1'b0;
      zz_rom_78[2] = 1'b0;
      zz_rom_78[3] = 1'b0;
      zz_rom_78[4] = 1'b0;
      zz_rom_78[5] = 1'b0;
      zz_rom_78[6] = 1'b0;
      zz_rom_78[7] = 1'b0;
      zz_rom_78[8] = 1'b0;
      zz_rom_78[9] = 1'b1;
      zz_rom_78[10] = 1'b1;
      zz_rom_78[11] = 1'b1;
      zz_rom_78[12] = 1'b1;
      zz_rom_78[13] = 1'b1;
      zz_rom_78[14] = 1'b1;
      zz_rom_78[15] = 1'b1;
      zz_rom_78[16] = 1'b1;
      zz_rom_78[17] = 1'b1;
      zz_rom_78[18] = 1'b1;
      zz_rom_78[19] = 1'b1;
      zz_rom_78[20] = 1'b1;
      zz_rom_78[21] = 1'b1;
      zz_rom_78[22] = 1'b1;
      zz_rom_78[23] = 1'b1;
      zz_rom_78[24] = 1'b1;
      zz_rom_78[25] = 1'b1;
      zz_rom_78[26] = 1'b1;
      zz_rom_78[27] = 1'b1;
      zz_rom_78[28] = 1'b1;
      zz_rom_78[29] = 1'b1;
      zz_rom_78[30] = 1'b1;
      zz_rom_78[31] = 1'b1;
      zz_rom_78[32] = 1'b1;
      zz_rom_78[33] = 1'b1;
      zz_rom_78[34] = 1'b1;
      zz_rom_78[35] = 1'b1;
      zz_rom_78[36] = 1'b1;
      zz_rom_78[37] = 1'b1;
      zz_rom_78[38] = 1'b1;
      zz_rom_78[39] = 1'b1;
      zz_rom_78[40] = 1'b1;
      zz_rom_78[41] = 1'b1;
      zz_rom_78[42] = 1'b1;
      zz_rom_78[43] = 1'b1;
      zz_rom_78[44] = 1'b1;
      zz_rom_78[45] = 1'b1;
      zz_rom_78[46] = 1'b1;
      zz_rom_78[47] = 1'b1;
      zz_rom_78[48] = 1'b1;
      zz_rom_78[49] = 1'b1;
      zz_rom_78[50] = 1'b1;
      zz_rom_78[51] = 1'b1;
      zz_rom_78[52] = 1'b1;
      zz_rom_78[53] = 1'b1;
      zz_rom_78[54] = 1'b1;
      zz_rom_78[55] = 1'b1;
      zz_rom_78[56] = 1'b1;
      zz_rom_78[57] = 1'b1;
      zz_rom_78[58] = 1'b1;
      zz_rom_78[59] = 1'b1;
      zz_rom_78[60] = 1'b1;
      zz_rom_78[61] = 1'b1;
      zz_rom_78[62] = 1'b1;
      zz_rom_78[63] = 1'b1;
      zz_rom_78[64] = 1'b1;
      zz_rom_78[65] = 1'b1;
      zz_rom_78[66] = 1'b1;
      zz_rom_78[67] = 1'b1;
      zz_rom_78[68] = 1'b1;
      zz_rom_78[69] = 1'b1;
      zz_rom_78[70] = 1'b1;
      zz_rom_78[71] = 1'b1;
      zz_rom_78[72] = 1'b1;
      zz_rom_78[73] = 1'b1;
      zz_rom_78[74] = 1'b1;
      zz_rom_78[75] = 1'b1;
      zz_rom_78[76] = 1'b1;
      zz_rom_78[77] = 1'b1;
      zz_rom_78[78] = 1'b1;
      zz_rom_78[79] = 1'b1;
      zz_rom_78[80] = 1'b1;
      zz_rom_78[81] = 1'b1;
      zz_rom_78[82] = 1'b1;
      zz_rom_78[83] = 1'b1;
      zz_rom_78[84] = 1'b1;
      zz_rom_78[85] = 1'b1;
      zz_rom_78[86] = 1'b1;
      zz_rom_78[87] = 1'b1;
      zz_rom_78[88] = 1'b1;
      zz_rom_78[89] = 1'b1;
      zz_rom_78[90] = 1'b1;
      zz_rom_78[91] = 1'b1;
      zz_rom_78[92] = 1'b0;
      zz_rom_78[93] = 1'b0;
      zz_rom_78[94] = 1'b0;
      zz_rom_78[95] = 1'b0;
      zz_rom_78[96] = 1'b0;
      zz_rom_78[97] = 1'b0;
      zz_rom_78[98] = 1'b0;
      zz_rom_78[99] = 1'b0;
    end
  endfunction
  wire [99:0] _zz_79;
  function [99:0] zz_rom_79(input dummy);
    begin
      zz_rom_79[0] = 1'b0;
      zz_rom_79[1] = 1'b0;
      zz_rom_79[2] = 1'b0;
      zz_rom_79[3] = 1'b0;
      zz_rom_79[4] = 1'b0;
      zz_rom_79[5] = 1'b0;
      zz_rom_79[6] = 1'b0;
      zz_rom_79[7] = 1'b0;
      zz_rom_79[8] = 1'b0;
      zz_rom_79[9] = 1'b0;
      zz_rom_79[10] = 1'b1;
      zz_rom_79[11] = 1'b1;
      zz_rom_79[12] = 1'b1;
      zz_rom_79[13] = 1'b1;
      zz_rom_79[14] = 1'b1;
      zz_rom_79[15] = 1'b1;
      zz_rom_79[16] = 1'b1;
      zz_rom_79[17] = 1'b1;
      zz_rom_79[18] = 1'b1;
      zz_rom_79[19] = 1'b1;
      zz_rom_79[20] = 1'b1;
      zz_rom_79[21] = 1'b1;
      zz_rom_79[22] = 1'b1;
      zz_rom_79[23] = 1'b1;
      zz_rom_79[24] = 1'b1;
      zz_rom_79[25] = 1'b1;
      zz_rom_79[26] = 1'b1;
      zz_rom_79[27] = 1'b1;
      zz_rom_79[28] = 1'b1;
      zz_rom_79[29] = 1'b1;
      zz_rom_79[30] = 1'b1;
      zz_rom_79[31] = 1'b1;
      zz_rom_79[32] = 1'b1;
      zz_rom_79[33] = 1'b1;
      zz_rom_79[34] = 1'b1;
      zz_rom_79[35] = 1'b1;
      zz_rom_79[36] = 1'b1;
      zz_rom_79[37] = 1'b1;
      zz_rom_79[38] = 1'b1;
      zz_rom_79[39] = 1'b1;
      zz_rom_79[40] = 1'b1;
      zz_rom_79[41] = 1'b1;
      zz_rom_79[42] = 1'b1;
      zz_rom_79[43] = 1'b1;
      zz_rom_79[44] = 1'b1;
      zz_rom_79[45] = 1'b1;
      zz_rom_79[46] = 1'b1;
      zz_rom_79[47] = 1'b1;
      zz_rom_79[48] = 1'b1;
      zz_rom_79[49] = 1'b1;
      zz_rom_79[50] = 1'b1;
      zz_rom_79[51] = 1'b1;
      zz_rom_79[52] = 1'b1;
      zz_rom_79[53] = 1'b1;
      zz_rom_79[54] = 1'b1;
      zz_rom_79[55] = 1'b1;
      zz_rom_79[56] = 1'b1;
      zz_rom_79[57] = 1'b1;
      zz_rom_79[58] = 1'b1;
      zz_rom_79[59] = 1'b1;
      zz_rom_79[60] = 1'b1;
      zz_rom_79[61] = 1'b1;
      zz_rom_79[62] = 1'b1;
      zz_rom_79[63] = 1'b1;
      zz_rom_79[64] = 1'b1;
      zz_rom_79[65] = 1'b1;
      zz_rom_79[66] = 1'b1;
      zz_rom_79[67] = 1'b1;
      zz_rom_79[68] = 1'b1;
      zz_rom_79[69] = 1'b1;
      zz_rom_79[70] = 1'b1;
      zz_rom_79[71] = 1'b1;
      zz_rom_79[72] = 1'b1;
      zz_rom_79[73] = 1'b1;
      zz_rom_79[74] = 1'b1;
      zz_rom_79[75] = 1'b1;
      zz_rom_79[76] = 1'b1;
      zz_rom_79[77] = 1'b1;
      zz_rom_79[78] = 1'b1;
      zz_rom_79[79] = 1'b1;
      zz_rom_79[80] = 1'b1;
      zz_rom_79[81] = 1'b1;
      zz_rom_79[82] = 1'b1;
      zz_rom_79[83] = 1'b1;
      zz_rom_79[84] = 1'b1;
      zz_rom_79[85] = 1'b1;
      zz_rom_79[86] = 1'b1;
      zz_rom_79[87] = 1'b1;
      zz_rom_79[88] = 1'b1;
      zz_rom_79[89] = 1'b1;
      zz_rom_79[90] = 1'b1;
      zz_rom_79[91] = 1'b0;
      zz_rom_79[92] = 1'b0;
      zz_rom_79[93] = 1'b0;
      zz_rom_79[94] = 1'b0;
      zz_rom_79[95] = 1'b0;
      zz_rom_79[96] = 1'b0;
      zz_rom_79[97] = 1'b0;
      zz_rom_79[98] = 1'b0;
      zz_rom_79[99] = 1'b0;
    end
  endfunction
  wire [99:0] _zz_80;
  function [99:0] zz_rom_80(input dummy);
    begin
      zz_rom_80[0] = 1'b0;
      zz_rom_80[1] = 1'b0;
      zz_rom_80[2] = 1'b0;
      zz_rom_80[3] = 1'b0;
      zz_rom_80[4] = 1'b0;
      zz_rom_80[5] = 1'b0;
      zz_rom_80[6] = 1'b0;
      zz_rom_80[7] = 1'b0;
      zz_rom_80[8] = 1'b0;
      zz_rom_80[9] = 1'b0;
      zz_rom_80[10] = 1'b1;
      zz_rom_80[11] = 1'b1;
      zz_rom_80[12] = 1'b1;
      zz_rom_80[13] = 1'b1;
      zz_rom_80[14] = 1'b1;
      zz_rom_80[15] = 1'b1;
      zz_rom_80[16] = 1'b1;
      zz_rom_80[17] = 1'b1;
      zz_rom_80[18] = 1'b1;
      zz_rom_80[19] = 1'b1;
      zz_rom_80[20] = 1'b1;
      zz_rom_80[21] = 1'b1;
      zz_rom_80[22] = 1'b1;
      zz_rom_80[23] = 1'b1;
      zz_rom_80[24] = 1'b1;
      zz_rom_80[25] = 1'b1;
      zz_rom_80[26] = 1'b1;
      zz_rom_80[27] = 1'b1;
      zz_rom_80[28] = 1'b1;
      zz_rom_80[29] = 1'b1;
      zz_rom_80[30] = 1'b1;
      zz_rom_80[31] = 1'b1;
      zz_rom_80[32] = 1'b1;
      zz_rom_80[33] = 1'b1;
      zz_rom_80[34] = 1'b1;
      zz_rom_80[35] = 1'b1;
      zz_rom_80[36] = 1'b1;
      zz_rom_80[37] = 1'b1;
      zz_rom_80[38] = 1'b1;
      zz_rom_80[39] = 1'b1;
      zz_rom_80[40] = 1'b1;
      zz_rom_80[41] = 1'b1;
      zz_rom_80[42] = 1'b1;
      zz_rom_80[43] = 1'b1;
      zz_rom_80[44] = 1'b1;
      zz_rom_80[45] = 1'b1;
      zz_rom_80[46] = 1'b1;
      zz_rom_80[47] = 1'b1;
      zz_rom_80[48] = 1'b1;
      zz_rom_80[49] = 1'b1;
      zz_rom_80[50] = 1'b1;
      zz_rom_80[51] = 1'b1;
      zz_rom_80[52] = 1'b1;
      zz_rom_80[53] = 1'b1;
      zz_rom_80[54] = 1'b1;
      zz_rom_80[55] = 1'b1;
      zz_rom_80[56] = 1'b1;
      zz_rom_80[57] = 1'b1;
      zz_rom_80[58] = 1'b1;
      zz_rom_80[59] = 1'b1;
      zz_rom_80[60] = 1'b1;
      zz_rom_80[61] = 1'b1;
      zz_rom_80[62] = 1'b1;
      zz_rom_80[63] = 1'b1;
      zz_rom_80[64] = 1'b1;
      zz_rom_80[65] = 1'b1;
      zz_rom_80[66] = 1'b1;
      zz_rom_80[67] = 1'b1;
      zz_rom_80[68] = 1'b1;
      zz_rom_80[69] = 1'b1;
      zz_rom_80[70] = 1'b1;
      zz_rom_80[71] = 1'b1;
      zz_rom_80[72] = 1'b1;
      zz_rom_80[73] = 1'b1;
      zz_rom_80[74] = 1'b1;
      zz_rom_80[75] = 1'b1;
      zz_rom_80[76] = 1'b1;
      zz_rom_80[77] = 1'b1;
      zz_rom_80[78] = 1'b1;
      zz_rom_80[79] = 1'b1;
      zz_rom_80[80] = 1'b1;
      zz_rom_80[81] = 1'b1;
      zz_rom_80[82] = 1'b1;
      zz_rom_80[83] = 1'b1;
      zz_rom_80[84] = 1'b1;
      zz_rom_80[85] = 1'b1;
      zz_rom_80[86] = 1'b1;
      zz_rom_80[87] = 1'b1;
      zz_rom_80[88] = 1'b1;
      zz_rom_80[89] = 1'b1;
      zz_rom_80[90] = 1'b1;
      zz_rom_80[91] = 1'b0;
      zz_rom_80[92] = 1'b0;
      zz_rom_80[93] = 1'b0;
      zz_rom_80[94] = 1'b0;
      zz_rom_80[95] = 1'b0;
      zz_rom_80[96] = 1'b0;
      zz_rom_80[97] = 1'b0;
      zz_rom_80[98] = 1'b0;
      zz_rom_80[99] = 1'b0;
    end
  endfunction
  wire [99:0] _zz_81;
  function [99:0] zz_rom_81(input dummy);
    begin
      zz_rom_81[0] = 1'b0;
      zz_rom_81[1] = 1'b0;
      zz_rom_81[2] = 1'b0;
      zz_rom_81[3] = 1'b0;
      zz_rom_81[4] = 1'b0;
      zz_rom_81[5] = 1'b0;
      zz_rom_81[6] = 1'b0;
      zz_rom_81[7] = 1'b0;
      zz_rom_81[8] = 1'b0;
      zz_rom_81[9] = 1'b0;
      zz_rom_81[10] = 1'b0;
      zz_rom_81[11] = 1'b1;
      zz_rom_81[12] = 1'b1;
      zz_rom_81[13] = 1'b1;
      zz_rom_81[14] = 1'b1;
      zz_rom_81[15] = 1'b1;
      zz_rom_81[16] = 1'b1;
      zz_rom_81[17] = 1'b1;
      zz_rom_81[18] = 1'b1;
      zz_rom_81[19] = 1'b1;
      zz_rom_81[20] = 1'b1;
      zz_rom_81[21] = 1'b1;
      zz_rom_81[22] = 1'b1;
      zz_rom_81[23] = 1'b1;
      zz_rom_81[24] = 1'b1;
      zz_rom_81[25] = 1'b1;
      zz_rom_81[26] = 1'b1;
      zz_rom_81[27] = 1'b1;
      zz_rom_81[28] = 1'b1;
      zz_rom_81[29] = 1'b1;
      zz_rom_81[30] = 1'b1;
      zz_rom_81[31] = 1'b1;
      zz_rom_81[32] = 1'b1;
      zz_rom_81[33] = 1'b1;
      zz_rom_81[34] = 1'b1;
      zz_rom_81[35] = 1'b1;
      zz_rom_81[36] = 1'b1;
      zz_rom_81[37] = 1'b1;
      zz_rom_81[38] = 1'b1;
      zz_rom_81[39] = 1'b1;
      zz_rom_81[40] = 1'b1;
      zz_rom_81[41] = 1'b1;
      zz_rom_81[42] = 1'b1;
      zz_rom_81[43] = 1'b1;
      zz_rom_81[44] = 1'b1;
      zz_rom_81[45] = 1'b1;
      zz_rom_81[46] = 1'b1;
      zz_rom_81[47] = 1'b1;
      zz_rom_81[48] = 1'b1;
      zz_rom_81[49] = 1'b1;
      zz_rom_81[50] = 1'b1;
      zz_rom_81[51] = 1'b1;
      zz_rom_81[52] = 1'b1;
      zz_rom_81[53] = 1'b1;
      zz_rom_81[54] = 1'b1;
      zz_rom_81[55] = 1'b1;
      zz_rom_81[56] = 1'b1;
      zz_rom_81[57] = 1'b1;
      zz_rom_81[58] = 1'b1;
      zz_rom_81[59] = 1'b1;
      zz_rom_81[60] = 1'b1;
      zz_rom_81[61] = 1'b1;
      zz_rom_81[62] = 1'b1;
      zz_rom_81[63] = 1'b1;
      zz_rom_81[64] = 1'b1;
      zz_rom_81[65] = 1'b1;
      zz_rom_81[66] = 1'b1;
      zz_rom_81[67] = 1'b1;
      zz_rom_81[68] = 1'b1;
      zz_rom_81[69] = 1'b1;
      zz_rom_81[70] = 1'b1;
      zz_rom_81[71] = 1'b1;
      zz_rom_81[72] = 1'b1;
      zz_rom_81[73] = 1'b1;
      zz_rom_81[74] = 1'b1;
      zz_rom_81[75] = 1'b1;
      zz_rom_81[76] = 1'b1;
      zz_rom_81[77] = 1'b1;
      zz_rom_81[78] = 1'b1;
      zz_rom_81[79] = 1'b1;
      zz_rom_81[80] = 1'b1;
      zz_rom_81[81] = 1'b1;
      zz_rom_81[82] = 1'b1;
      zz_rom_81[83] = 1'b1;
      zz_rom_81[84] = 1'b1;
      zz_rom_81[85] = 1'b1;
      zz_rom_81[86] = 1'b1;
      zz_rom_81[87] = 1'b1;
      zz_rom_81[88] = 1'b1;
      zz_rom_81[89] = 1'b1;
      zz_rom_81[90] = 1'b0;
      zz_rom_81[91] = 1'b0;
      zz_rom_81[92] = 1'b0;
      zz_rom_81[93] = 1'b0;
      zz_rom_81[94] = 1'b0;
      zz_rom_81[95] = 1'b0;
      zz_rom_81[96] = 1'b0;
      zz_rom_81[97] = 1'b0;
      zz_rom_81[98] = 1'b0;
      zz_rom_81[99] = 1'b0;
    end
  endfunction
  wire [99:0] _zz_82;
  function [99:0] zz_rom_82(input dummy);
    begin
      zz_rom_82[0] = 1'b0;
      zz_rom_82[1] = 1'b0;
      zz_rom_82[2] = 1'b0;
      zz_rom_82[3] = 1'b0;
      zz_rom_82[4] = 1'b0;
      zz_rom_82[5] = 1'b0;
      zz_rom_82[6] = 1'b0;
      zz_rom_82[7] = 1'b0;
      zz_rom_82[8] = 1'b0;
      zz_rom_82[9] = 1'b0;
      zz_rom_82[10] = 1'b0;
      zz_rom_82[11] = 1'b0;
      zz_rom_82[12] = 1'b1;
      zz_rom_82[13] = 1'b1;
      zz_rom_82[14] = 1'b1;
      zz_rom_82[15] = 1'b1;
      zz_rom_82[16] = 1'b1;
      zz_rom_82[17] = 1'b1;
      zz_rom_82[18] = 1'b1;
      zz_rom_82[19] = 1'b1;
      zz_rom_82[20] = 1'b1;
      zz_rom_82[21] = 1'b1;
      zz_rom_82[22] = 1'b1;
      zz_rom_82[23] = 1'b1;
      zz_rom_82[24] = 1'b1;
      zz_rom_82[25] = 1'b1;
      zz_rom_82[26] = 1'b1;
      zz_rom_82[27] = 1'b1;
      zz_rom_82[28] = 1'b1;
      zz_rom_82[29] = 1'b1;
      zz_rom_82[30] = 1'b1;
      zz_rom_82[31] = 1'b1;
      zz_rom_82[32] = 1'b1;
      zz_rom_82[33] = 1'b1;
      zz_rom_82[34] = 1'b1;
      zz_rom_82[35] = 1'b1;
      zz_rom_82[36] = 1'b1;
      zz_rom_82[37] = 1'b1;
      zz_rom_82[38] = 1'b1;
      zz_rom_82[39] = 1'b1;
      zz_rom_82[40] = 1'b1;
      zz_rom_82[41] = 1'b1;
      zz_rom_82[42] = 1'b1;
      zz_rom_82[43] = 1'b1;
      zz_rom_82[44] = 1'b1;
      zz_rom_82[45] = 1'b1;
      zz_rom_82[46] = 1'b1;
      zz_rom_82[47] = 1'b1;
      zz_rom_82[48] = 1'b1;
      zz_rom_82[49] = 1'b1;
      zz_rom_82[50] = 1'b1;
      zz_rom_82[51] = 1'b1;
      zz_rom_82[52] = 1'b1;
      zz_rom_82[53] = 1'b1;
      zz_rom_82[54] = 1'b1;
      zz_rom_82[55] = 1'b1;
      zz_rom_82[56] = 1'b1;
      zz_rom_82[57] = 1'b1;
      zz_rom_82[58] = 1'b1;
      zz_rom_82[59] = 1'b1;
      zz_rom_82[60] = 1'b1;
      zz_rom_82[61] = 1'b1;
      zz_rom_82[62] = 1'b1;
      zz_rom_82[63] = 1'b1;
      zz_rom_82[64] = 1'b1;
      zz_rom_82[65] = 1'b1;
      zz_rom_82[66] = 1'b1;
      zz_rom_82[67] = 1'b1;
      zz_rom_82[68] = 1'b1;
      zz_rom_82[69] = 1'b1;
      zz_rom_82[70] = 1'b1;
      zz_rom_82[71] = 1'b1;
      zz_rom_82[72] = 1'b1;
      zz_rom_82[73] = 1'b1;
      zz_rom_82[74] = 1'b1;
      zz_rom_82[75] = 1'b1;
      zz_rom_82[76] = 1'b1;
      zz_rom_82[77] = 1'b1;
      zz_rom_82[78] = 1'b1;
      zz_rom_82[79] = 1'b1;
      zz_rom_82[80] = 1'b1;
      zz_rom_82[81] = 1'b1;
      zz_rom_82[82] = 1'b1;
      zz_rom_82[83] = 1'b1;
      zz_rom_82[84] = 1'b1;
      zz_rom_82[85] = 1'b1;
      zz_rom_82[86] = 1'b1;
      zz_rom_82[87] = 1'b1;
      zz_rom_82[88] = 1'b1;
      zz_rom_82[89] = 1'b0;
      zz_rom_82[90] = 1'b0;
      zz_rom_82[91] = 1'b0;
      zz_rom_82[92] = 1'b0;
      zz_rom_82[93] = 1'b0;
      zz_rom_82[94] = 1'b0;
      zz_rom_82[95] = 1'b0;
      zz_rom_82[96] = 1'b0;
      zz_rom_82[97] = 1'b0;
      zz_rom_82[98] = 1'b0;
      zz_rom_82[99] = 1'b0;
    end
  endfunction
  wire [99:0] _zz_83;
  function [99:0] zz_rom_83(input dummy);
    begin
      zz_rom_83[0] = 1'b0;
      zz_rom_83[1] = 1'b0;
      zz_rom_83[2] = 1'b0;
      zz_rom_83[3] = 1'b0;
      zz_rom_83[4] = 1'b0;
      zz_rom_83[5] = 1'b0;
      zz_rom_83[6] = 1'b0;
      zz_rom_83[7] = 1'b0;
      zz_rom_83[8] = 1'b0;
      zz_rom_83[9] = 1'b0;
      zz_rom_83[10] = 1'b0;
      zz_rom_83[11] = 1'b0;
      zz_rom_83[12] = 1'b0;
      zz_rom_83[13] = 1'b1;
      zz_rom_83[14] = 1'b1;
      zz_rom_83[15] = 1'b1;
      zz_rom_83[16] = 1'b1;
      zz_rom_83[17] = 1'b1;
      zz_rom_83[18] = 1'b1;
      zz_rom_83[19] = 1'b1;
      zz_rom_83[20] = 1'b1;
      zz_rom_83[21] = 1'b1;
      zz_rom_83[22] = 1'b1;
      zz_rom_83[23] = 1'b1;
      zz_rom_83[24] = 1'b1;
      zz_rom_83[25] = 1'b1;
      zz_rom_83[26] = 1'b1;
      zz_rom_83[27] = 1'b1;
      zz_rom_83[28] = 1'b1;
      zz_rom_83[29] = 1'b1;
      zz_rom_83[30] = 1'b1;
      zz_rom_83[31] = 1'b1;
      zz_rom_83[32] = 1'b1;
      zz_rom_83[33] = 1'b1;
      zz_rom_83[34] = 1'b1;
      zz_rom_83[35] = 1'b1;
      zz_rom_83[36] = 1'b1;
      zz_rom_83[37] = 1'b1;
      zz_rom_83[38] = 1'b1;
      zz_rom_83[39] = 1'b1;
      zz_rom_83[40] = 1'b1;
      zz_rom_83[41] = 1'b1;
      zz_rom_83[42] = 1'b1;
      zz_rom_83[43] = 1'b1;
      zz_rom_83[44] = 1'b1;
      zz_rom_83[45] = 1'b1;
      zz_rom_83[46] = 1'b1;
      zz_rom_83[47] = 1'b1;
      zz_rom_83[48] = 1'b1;
      zz_rom_83[49] = 1'b1;
      zz_rom_83[50] = 1'b1;
      zz_rom_83[51] = 1'b1;
      zz_rom_83[52] = 1'b1;
      zz_rom_83[53] = 1'b1;
      zz_rom_83[54] = 1'b1;
      zz_rom_83[55] = 1'b1;
      zz_rom_83[56] = 1'b1;
      zz_rom_83[57] = 1'b1;
      zz_rom_83[58] = 1'b1;
      zz_rom_83[59] = 1'b1;
      zz_rom_83[60] = 1'b1;
      zz_rom_83[61] = 1'b1;
      zz_rom_83[62] = 1'b1;
      zz_rom_83[63] = 1'b1;
      zz_rom_83[64] = 1'b1;
      zz_rom_83[65] = 1'b1;
      zz_rom_83[66] = 1'b1;
      zz_rom_83[67] = 1'b1;
      zz_rom_83[68] = 1'b1;
      zz_rom_83[69] = 1'b1;
      zz_rom_83[70] = 1'b1;
      zz_rom_83[71] = 1'b1;
      zz_rom_83[72] = 1'b1;
      zz_rom_83[73] = 1'b1;
      zz_rom_83[74] = 1'b1;
      zz_rom_83[75] = 1'b1;
      zz_rom_83[76] = 1'b1;
      zz_rom_83[77] = 1'b1;
      zz_rom_83[78] = 1'b1;
      zz_rom_83[79] = 1'b1;
      zz_rom_83[80] = 1'b1;
      zz_rom_83[81] = 1'b1;
      zz_rom_83[82] = 1'b1;
      zz_rom_83[83] = 1'b1;
      zz_rom_83[84] = 1'b1;
      zz_rom_83[85] = 1'b1;
      zz_rom_83[86] = 1'b1;
      zz_rom_83[87] = 1'b1;
      zz_rom_83[88] = 1'b0;
      zz_rom_83[89] = 1'b0;
      zz_rom_83[90] = 1'b0;
      zz_rom_83[91] = 1'b0;
      zz_rom_83[92] = 1'b0;
      zz_rom_83[93] = 1'b0;
      zz_rom_83[94] = 1'b0;
      zz_rom_83[95] = 1'b0;
      zz_rom_83[96] = 1'b0;
      zz_rom_83[97] = 1'b0;
      zz_rom_83[98] = 1'b0;
      zz_rom_83[99] = 1'b0;
    end
  endfunction
  wire [99:0] _zz_84;
  function [99:0] zz_rom_84(input dummy);
    begin
      zz_rom_84[0] = 1'b0;
      zz_rom_84[1] = 1'b0;
      zz_rom_84[2] = 1'b0;
      zz_rom_84[3] = 1'b0;
      zz_rom_84[4] = 1'b0;
      zz_rom_84[5] = 1'b0;
      zz_rom_84[6] = 1'b0;
      zz_rom_84[7] = 1'b0;
      zz_rom_84[8] = 1'b0;
      zz_rom_84[9] = 1'b0;
      zz_rom_84[10] = 1'b0;
      zz_rom_84[11] = 1'b0;
      zz_rom_84[12] = 1'b0;
      zz_rom_84[13] = 1'b0;
      zz_rom_84[14] = 1'b1;
      zz_rom_84[15] = 1'b1;
      zz_rom_84[16] = 1'b1;
      zz_rom_84[17] = 1'b1;
      zz_rom_84[18] = 1'b1;
      zz_rom_84[19] = 1'b1;
      zz_rom_84[20] = 1'b1;
      zz_rom_84[21] = 1'b1;
      zz_rom_84[22] = 1'b1;
      zz_rom_84[23] = 1'b1;
      zz_rom_84[24] = 1'b1;
      zz_rom_84[25] = 1'b1;
      zz_rom_84[26] = 1'b1;
      zz_rom_84[27] = 1'b1;
      zz_rom_84[28] = 1'b1;
      zz_rom_84[29] = 1'b1;
      zz_rom_84[30] = 1'b1;
      zz_rom_84[31] = 1'b1;
      zz_rom_84[32] = 1'b1;
      zz_rom_84[33] = 1'b1;
      zz_rom_84[34] = 1'b1;
      zz_rom_84[35] = 1'b1;
      zz_rom_84[36] = 1'b1;
      zz_rom_84[37] = 1'b1;
      zz_rom_84[38] = 1'b1;
      zz_rom_84[39] = 1'b1;
      zz_rom_84[40] = 1'b1;
      zz_rom_84[41] = 1'b1;
      zz_rom_84[42] = 1'b1;
      zz_rom_84[43] = 1'b1;
      zz_rom_84[44] = 1'b1;
      zz_rom_84[45] = 1'b1;
      zz_rom_84[46] = 1'b1;
      zz_rom_84[47] = 1'b1;
      zz_rom_84[48] = 1'b1;
      zz_rom_84[49] = 1'b1;
      zz_rom_84[50] = 1'b1;
      zz_rom_84[51] = 1'b1;
      zz_rom_84[52] = 1'b1;
      zz_rom_84[53] = 1'b1;
      zz_rom_84[54] = 1'b1;
      zz_rom_84[55] = 1'b1;
      zz_rom_84[56] = 1'b1;
      zz_rom_84[57] = 1'b1;
      zz_rom_84[58] = 1'b1;
      zz_rom_84[59] = 1'b1;
      zz_rom_84[60] = 1'b1;
      zz_rom_84[61] = 1'b1;
      zz_rom_84[62] = 1'b1;
      zz_rom_84[63] = 1'b1;
      zz_rom_84[64] = 1'b1;
      zz_rom_84[65] = 1'b1;
      zz_rom_84[66] = 1'b1;
      zz_rom_84[67] = 1'b1;
      zz_rom_84[68] = 1'b1;
      zz_rom_84[69] = 1'b1;
      zz_rom_84[70] = 1'b1;
      zz_rom_84[71] = 1'b1;
      zz_rom_84[72] = 1'b1;
      zz_rom_84[73] = 1'b1;
      zz_rom_84[74] = 1'b1;
      zz_rom_84[75] = 1'b1;
      zz_rom_84[76] = 1'b1;
      zz_rom_84[77] = 1'b1;
      zz_rom_84[78] = 1'b1;
      zz_rom_84[79] = 1'b1;
      zz_rom_84[80] = 1'b1;
      zz_rom_84[81] = 1'b1;
      zz_rom_84[82] = 1'b1;
      zz_rom_84[83] = 1'b1;
      zz_rom_84[84] = 1'b1;
      zz_rom_84[85] = 1'b1;
      zz_rom_84[86] = 1'b1;
      zz_rom_84[87] = 1'b0;
      zz_rom_84[88] = 1'b0;
      zz_rom_84[89] = 1'b0;
      zz_rom_84[90] = 1'b0;
      zz_rom_84[91] = 1'b0;
      zz_rom_84[92] = 1'b0;
      zz_rom_84[93] = 1'b0;
      zz_rom_84[94] = 1'b0;
      zz_rom_84[95] = 1'b0;
      zz_rom_84[96] = 1'b0;
      zz_rom_84[97] = 1'b0;
      zz_rom_84[98] = 1'b0;
      zz_rom_84[99] = 1'b0;
    end
  endfunction
  wire [99:0] _zz_85;
  function [99:0] zz_rom_85(input dummy);
    begin
      zz_rom_85[0] = 1'b0;
      zz_rom_85[1] = 1'b0;
      zz_rom_85[2] = 1'b0;
      zz_rom_85[3] = 1'b0;
      zz_rom_85[4] = 1'b0;
      zz_rom_85[5] = 1'b0;
      zz_rom_85[6] = 1'b0;
      zz_rom_85[7] = 1'b0;
      zz_rom_85[8] = 1'b0;
      zz_rom_85[9] = 1'b0;
      zz_rom_85[10] = 1'b0;
      zz_rom_85[11] = 1'b0;
      zz_rom_85[12] = 1'b0;
      zz_rom_85[13] = 1'b0;
      zz_rom_85[14] = 1'b0;
      zz_rom_85[15] = 1'b1;
      zz_rom_85[16] = 1'b1;
      zz_rom_85[17] = 1'b1;
      zz_rom_85[18] = 1'b1;
      zz_rom_85[19] = 1'b1;
      zz_rom_85[20] = 1'b1;
      zz_rom_85[21] = 1'b1;
      zz_rom_85[22] = 1'b1;
      zz_rom_85[23] = 1'b1;
      zz_rom_85[24] = 1'b1;
      zz_rom_85[25] = 1'b1;
      zz_rom_85[26] = 1'b1;
      zz_rom_85[27] = 1'b1;
      zz_rom_85[28] = 1'b1;
      zz_rom_85[29] = 1'b1;
      zz_rom_85[30] = 1'b1;
      zz_rom_85[31] = 1'b1;
      zz_rom_85[32] = 1'b1;
      zz_rom_85[33] = 1'b1;
      zz_rom_85[34] = 1'b1;
      zz_rom_85[35] = 1'b1;
      zz_rom_85[36] = 1'b1;
      zz_rom_85[37] = 1'b1;
      zz_rom_85[38] = 1'b1;
      zz_rom_85[39] = 1'b1;
      zz_rom_85[40] = 1'b1;
      zz_rom_85[41] = 1'b1;
      zz_rom_85[42] = 1'b1;
      zz_rom_85[43] = 1'b1;
      zz_rom_85[44] = 1'b1;
      zz_rom_85[45] = 1'b1;
      zz_rom_85[46] = 1'b1;
      zz_rom_85[47] = 1'b1;
      zz_rom_85[48] = 1'b1;
      zz_rom_85[49] = 1'b1;
      zz_rom_85[50] = 1'b1;
      zz_rom_85[51] = 1'b1;
      zz_rom_85[52] = 1'b1;
      zz_rom_85[53] = 1'b1;
      zz_rom_85[54] = 1'b1;
      zz_rom_85[55] = 1'b1;
      zz_rom_85[56] = 1'b1;
      zz_rom_85[57] = 1'b1;
      zz_rom_85[58] = 1'b1;
      zz_rom_85[59] = 1'b1;
      zz_rom_85[60] = 1'b1;
      zz_rom_85[61] = 1'b1;
      zz_rom_85[62] = 1'b1;
      zz_rom_85[63] = 1'b1;
      zz_rom_85[64] = 1'b1;
      zz_rom_85[65] = 1'b1;
      zz_rom_85[66] = 1'b1;
      zz_rom_85[67] = 1'b1;
      zz_rom_85[68] = 1'b1;
      zz_rom_85[69] = 1'b1;
      zz_rom_85[70] = 1'b1;
      zz_rom_85[71] = 1'b1;
      zz_rom_85[72] = 1'b1;
      zz_rom_85[73] = 1'b1;
      zz_rom_85[74] = 1'b1;
      zz_rom_85[75] = 1'b1;
      zz_rom_85[76] = 1'b1;
      zz_rom_85[77] = 1'b1;
      zz_rom_85[78] = 1'b1;
      zz_rom_85[79] = 1'b1;
      zz_rom_85[80] = 1'b1;
      zz_rom_85[81] = 1'b1;
      zz_rom_85[82] = 1'b1;
      zz_rom_85[83] = 1'b1;
      zz_rom_85[84] = 1'b1;
      zz_rom_85[85] = 1'b1;
      zz_rom_85[86] = 1'b0;
      zz_rom_85[87] = 1'b0;
      zz_rom_85[88] = 1'b0;
      zz_rom_85[89] = 1'b0;
      zz_rom_85[90] = 1'b0;
      zz_rom_85[91] = 1'b0;
      zz_rom_85[92] = 1'b0;
      zz_rom_85[93] = 1'b0;
      zz_rom_85[94] = 1'b0;
      zz_rom_85[95] = 1'b0;
      zz_rom_85[96] = 1'b0;
      zz_rom_85[97] = 1'b0;
      zz_rom_85[98] = 1'b0;
      zz_rom_85[99] = 1'b0;
    end
  endfunction
  wire [99:0] _zz_86;
  function [99:0] zz_rom_86(input dummy);
    begin
      zz_rom_86[0] = 1'b0;
      zz_rom_86[1] = 1'b0;
      zz_rom_86[2] = 1'b0;
      zz_rom_86[3] = 1'b0;
      zz_rom_86[4] = 1'b0;
      zz_rom_86[5] = 1'b0;
      zz_rom_86[6] = 1'b0;
      zz_rom_86[7] = 1'b0;
      zz_rom_86[8] = 1'b0;
      zz_rom_86[9] = 1'b0;
      zz_rom_86[10] = 1'b0;
      zz_rom_86[11] = 1'b0;
      zz_rom_86[12] = 1'b0;
      zz_rom_86[13] = 1'b0;
      zz_rom_86[14] = 1'b0;
      zz_rom_86[15] = 1'b0;
      zz_rom_86[16] = 1'b1;
      zz_rom_86[17] = 1'b1;
      zz_rom_86[18] = 1'b1;
      zz_rom_86[19] = 1'b1;
      zz_rom_86[20] = 1'b1;
      zz_rom_86[21] = 1'b1;
      zz_rom_86[22] = 1'b1;
      zz_rom_86[23] = 1'b1;
      zz_rom_86[24] = 1'b1;
      zz_rom_86[25] = 1'b1;
      zz_rom_86[26] = 1'b1;
      zz_rom_86[27] = 1'b1;
      zz_rom_86[28] = 1'b1;
      zz_rom_86[29] = 1'b1;
      zz_rom_86[30] = 1'b1;
      zz_rom_86[31] = 1'b1;
      zz_rom_86[32] = 1'b1;
      zz_rom_86[33] = 1'b1;
      zz_rom_86[34] = 1'b1;
      zz_rom_86[35] = 1'b1;
      zz_rom_86[36] = 1'b1;
      zz_rom_86[37] = 1'b1;
      zz_rom_86[38] = 1'b1;
      zz_rom_86[39] = 1'b1;
      zz_rom_86[40] = 1'b1;
      zz_rom_86[41] = 1'b1;
      zz_rom_86[42] = 1'b1;
      zz_rom_86[43] = 1'b1;
      zz_rom_86[44] = 1'b1;
      zz_rom_86[45] = 1'b1;
      zz_rom_86[46] = 1'b1;
      zz_rom_86[47] = 1'b1;
      zz_rom_86[48] = 1'b1;
      zz_rom_86[49] = 1'b1;
      zz_rom_86[50] = 1'b1;
      zz_rom_86[51] = 1'b1;
      zz_rom_86[52] = 1'b1;
      zz_rom_86[53] = 1'b1;
      zz_rom_86[54] = 1'b1;
      zz_rom_86[55] = 1'b1;
      zz_rom_86[56] = 1'b1;
      zz_rom_86[57] = 1'b1;
      zz_rom_86[58] = 1'b1;
      zz_rom_86[59] = 1'b1;
      zz_rom_86[60] = 1'b1;
      zz_rom_86[61] = 1'b1;
      zz_rom_86[62] = 1'b1;
      zz_rom_86[63] = 1'b1;
      zz_rom_86[64] = 1'b1;
      zz_rom_86[65] = 1'b1;
      zz_rom_86[66] = 1'b1;
      zz_rom_86[67] = 1'b1;
      zz_rom_86[68] = 1'b1;
      zz_rom_86[69] = 1'b1;
      zz_rom_86[70] = 1'b1;
      zz_rom_86[71] = 1'b1;
      zz_rom_86[72] = 1'b1;
      zz_rom_86[73] = 1'b1;
      zz_rom_86[74] = 1'b1;
      zz_rom_86[75] = 1'b1;
      zz_rom_86[76] = 1'b1;
      zz_rom_86[77] = 1'b1;
      zz_rom_86[78] = 1'b1;
      zz_rom_86[79] = 1'b1;
      zz_rom_86[80] = 1'b1;
      zz_rom_86[81] = 1'b1;
      zz_rom_86[82] = 1'b1;
      zz_rom_86[83] = 1'b1;
      zz_rom_86[84] = 1'b1;
      zz_rom_86[85] = 1'b0;
      zz_rom_86[86] = 1'b0;
      zz_rom_86[87] = 1'b0;
      zz_rom_86[88] = 1'b0;
      zz_rom_86[89] = 1'b0;
      zz_rom_86[90] = 1'b0;
      zz_rom_86[91] = 1'b0;
      zz_rom_86[92] = 1'b0;
      zz_rom_86[93] = 1'b0;
      zz_rom_86[94] = 1'b0;
      zz_rom_86[95] = 1'b0;
      zz_rom_86[96] = 1'b0;
      zz_rom_86[97] = 1'b0;
      zz_rom_86[98] = 1'b0;
      zz_rom_86[99] = 1'b0;
    end
  endfunction
  wire [99:0] _zz_87;
  function [99:0] zz_rom_87(input dummy);
    begin
      zz_rom_87[0] = 1'b0;
      zz_rom_87[1] = 1'b0;
      zz_rom_87[2] = 1'b0;
      zz_rom_87[3] = 1'b0;
      zz_rom_87[4] = 1'b0;
      zz_rom_87[5] = 1'b0;
      zz_rom_87[6] = 1'b0;
      zz_rom_87[7] = 1'b0;
      zz_rom_87[8] = 1'b0;
      zz_rom_87[9] = 1'b0;
      zz_rom_87[10] = 1'b0;
      zz_rom_87[11] = 1'b0;
      zz_rom_87[12] = 1'b0;
      zz_rom_87[13] = 1'b0;
      zz_rom_87[14] = 1'b0;
      zz_rom_87[15] = 1'b0;
      zz_rom_87[16] = 1'b0;
      zz_rom_87[17] = 1'b1;
      zz_rom_87[18] = 1'b1;
      zz_rom_87[19] = 1'b1;
      zz_rom_87[20] = 1'b1;
      zz_rom_87[21] = 1'b1;
      zz_rom_87[22] = 1'b1;
      zz_rom_87[23] = 1'b1;
      zz_rom_87[24] = 1'b1;
      zz_rom_87[25] = 1'b1;
      zz_rom_87[26] = 1'b1;
      zz_rom_87[27] = 1'b1;
      zz_rom_87[28] = 1'b1;
      zz_rom_87[29] = 1'b1;
      zz_rom_87[30] = 1'b1;
      zz_rom_87[31] = 1'b1;
      zz_rom_87[32] = 1'b1;
      zz_rom_87[33] = 1'b1;
      zz_rom_87[34] = 1'b1;
      zz_rom_87[35] = 1'b1;
      zz_rom_87[36] = 1'b1;
      zz_rom_87[37] = 1'b1;
      zz_rom_87[38] = 1'b1;
      zz_rom_87[39] = 1'b1;
      zz_rom_87[40] = 1'b1;
      zz_rom_87[41] = 1'b1;
      zz_rom_87[42] = 1'b1;
      zz_rom_87[43] = 1'b1;
      zz_rom_87[44] = 1'b1;
      zz_rom_87[45] = 1'b1;
      zz_rom_87[46] = 1'b1;
      zz_rom_87[47] = 1'b1;
      zz_rom_87[48] = 1'b1;
      zz_rom_87[49] = 1'b1;
      zz_rom_87[50] = 1'b1;
      zz_rom_87[51] = 1'b1;
      zz_rom_87[52] = 1'b1;
      zz_rom_87[53] = 1'b1;
      zz_rom_87[54] = 1'b1;
      zz_rom_87[55] = 1'b1;
      zz_rom_87[56] = 1'b1;
      zz_rom_87[57] = 1'b1;
      zz_rom_87[58] = 1'b1;
      zz_rom_87[59] = 1'b1;
      zz_rom_87[60] = 1'b1;
      zz_rom_87[61] = 1'b1;
      zz_rom_87[62] = 1'b1;
      zz_rom_87[63] = 1'b1;
      zz_rom_87[64] = 1'b1;
      zz_rom_87[65] = 1'b1;
      zz_rom_87[66] = 1'b1;
      zz_rom_87[67] = 1'b1;
      zz_rom_87[68] = 1'b1;
      zz_rom_87[69] = 1'b1;
      zz_rom_87[70] = 1'b1;
      zz_rom_87[71] = 1'b1;
      zz_rom_87[72] = 1'b1;
      zz_rom_87[73] = 1'b1;
      zz_rom_87[74] = 1'b1;
      zz_rom_87[75] = 1'b1;
      zz_rom_87[76] = 1'b1;
      zz_rom_87[77] = 1'b1;
      zz_rom_87[78] = 1'b1;
      zz_rom_87[79] = 1'b1;
      zz_rom_87[80] = 1'b1;
      zz_rom_87[81] = 1'b1;
      zz_rom_87[82] = 1'b1;
      zz_rom_87[83] = 1'b1;
      zz_rom_87[84] = 1'b0;
      zz_rom_87[85] = 1'b0;
      zz_rom_87[86] = 1'b0;
      zz_rom_87[87] = 1'b0;
      zz_rom_87[88] = 1'b0;
      zz_rom_87[89] = 1'b0;
      zz_rom_87[90] = 1'b0;
      zz_rom_87[91] = 1'b0;
      zz_rom_87[92] = 1'b0;
      zz_rom_87[93] = 1'b0;
      zz_rom_87[94] = 1'b0;
      zz_rom_87[95] = 1'b0;
      zz_rom_87[96] = 1'b0;
      zz_rom_87[97] = 1'b0;
      zz_rom_87[98] = 1'b0;
      zz_rom_87[99] = 1'b0;
    end
  endfunction
  wire [99:0] _zz_88;
  function [99:0] zz_rom_88(input dummy);
    begin
      zz_rom_88[0] = 1'b0;
      zz_rom_88[1] = 1'b0;
      zz_rom_88[2] = 1'b0;
      zz_rom_88[3] = 1'b0;
      zz_rom_88[4] = 1'b0;
      zz_rom_88[5] = 1'b0;
      zz_rom_88[6] = 1'b0;
      zz_rom_88[7] = 1'b0;
      zz_rom_88[8] = 1'b0;
      zz_rom_88[9] = 1'b0;
      zz_rom_88[10] = 1'b0;
      zz_rom_88[11] = 1'b0;
      zz_rom_88[12] = 1'b0;
      zz_rom_88[13] = 1'b0;
      zz_rom_88[14] = 1'b0;
      zz_rom_88[15] = 1'b0;
      zz_rom_88[16] = 1'b0;
      zz_rom_88[17] = 1'b0;
      zz_rom_88[18] = 1'b1;
      zz_rom_88[19] = 1'b1;
      zz_rom_88[20] = 1'b1;
      zz_rom_88[21] = 1'b1;
      zz_rom_88[22] = 1'b1;
      zz_rom_88[23] = 1'b1;
      zz_rom_88[24] = 1'b1;
      zz_rom_88[25] = 1'b1;
      zz_rom_88[26] = 1'b1;
      zz_rom_88[27] = 1'b1;
      zz_rom_88[28] = 1'b1;
      zz_rom_88[29] = 1'b1;
      zz_rom_88[30] = 1'b1;
      zz_rom_88[31] = 1'b1;
      zz_rom_88[32] = 1'b1;
      zz_rom_88[33] = 1'b1;
      zz_rom_88[34] = 1'b1;
      zz_rom_88[35] = 1'b1;
      zz_rom_88[36] = 1'b1;
      zz_rom_88[37] = 1'b1;
      zz_rom_88[38] = 1'b1;
      zz_rom_88[39] = 1'b1;
      zz_rom_88[40] = 1'b1;
      zz_rom_88[41] = 1'b1;
      zz_rom_88[42] = 1'b1;
      zz_rom_88[43] = 1'b1;
      zz_rom_88[44] = 1'b1;
      zz_rom_88[45] = 1'b1;
      zz_rom_88[46] = 1'b1;
      zz_rom_88[47] = 1'b1;
      zz_rom_88[48] = 1'b1;
      zz_rom_88[49] = 1'b1;
      zz_rom_88[50] = 1'b1;
      zz_rom_88[51] = 1'b1;
      zz_rom_88[52] = 1'b1;
      zz_rom_88[53] = 1'b1;
      zz_rom_88[54] = 1'b1;
      zz_rom_88[55] = 1'b1;
      zz_rom_88[56] = 1'b1;
      zz_rom_88[57] = 1'b1;
      zz_rom_88[58] = 1'b1;
      zz_rom_88[59] = 1'b1;
      zz_rom_88[60] = 1'b1;
      zz_rom_88[61] = 1'b1;
      zz_rom_88[62] = 1'b1;
      zz_rom_88[63] = 1'b1;
      zz_rom_88[64] = 1'b1;
      zz_rom_88[65] = 1'b1;
      zz_rom_88[66] = 1'b1;
      zz_rom_88[67] = 1'b1;
      zz_rom_88[68] = 1'b1;
      zz_rom_88[69] = 1'b1;
      zz_rom_88[70] = 1'b1;
      zz_rom_88[71] = 1'b1;
      zz_rom_88[72] = 1'b1;
      zz_rom_88[73] = 1'b1;
      zz_rom_88[74] = 1'b1;
      zz_rom_88[75] = 1'b1;
      zz_rom_88[76] = 1'b1;
      zz_rom_88[77] = 1'b1;
      zz_rom_88[78] = 1'b1;
      zz_rom_88[79] = 1'b1;
      zz_rom_88[80] = 1'b1;
      zz_rom_88[81] = 1'b1;
      zz_rom_88[82] = 1'b1;
      zz_rom_88[83] = 1'b0;
      zz_rom_88[84] = 1'b0;
      zz_rom_88[85] = 1'b0;
      zz_rom_88[86] = 1'b0;
      zz_rom_88[87] = 1'b0;
      zz_rom_88[88] = 1'b0;
      zz_rom_88[89] = 1'b0;
      zz_rom_88[90] = 1'b0;
      zz_rom_88[91] = 1'b0;
      zz_rom_88[92] = 1'b0;
      zz_rom_88[93] = 1'b0;
      zz_rom_88[94] = 1'b0;
      zz_rom_88[95] = 1'b0;
      zz_rom_88[96] = 1'b0;
      zz_rom_88[97] = 1'b0;
      zz_rom_88[98] = 1'b0;
      zz_rom_88[99] = 1'b0;
    end
  endfunction
  wire [99:0] _zz_89;
  function [99:0] zz_rom_89(input dummy);
    begin
      zz_rom_89[0] = 1'b0;
      zz_rom_89[1] = 1'b0;
      zz_rom_89[2] = 1'b0;
      zz_rom_89[3] = 1'b0;
      zz_rom_89[4] = 1'b0;
      zz_rom_89[5] = 1'b0;
      zz_rom_89[6] = 1'b0;
      zz_rom_89[7] = 1'b0;
      zz_rom_89[8] = 1'b0;
      zz_rom_89[9] = 1'b0;
      zz_rom_89[10] = 1'b0;
      zz_rom_89[11] = 1'b0;
      zz_rom_89[12] = 1'b0;
      zz_rom_89[13] = 1'b0;
      zz_rom_89[14] = 1'b0;
      zz_rom_89[15] = 1'b0;
      zz_rom_89[16] = 1'b0;
      zz_rom_89[17] = 1'b0;
      zz_rom_89[18] = 1'b0;
      zz_rom_89[19] = 1'b1;
      zz_rom_89[20] = 1'b1;
      zz_rom_89[21] = 1'b1;
      zz_rom_89[22] = 1'b1;
      zz_rom_89[23] = 1'b1;
      zz_rom_89[24] = 1'b1;
      zz_rom_89[25] = 1'b1;
      zz_rom_89[26] = 1'b1;
      zz_rom_89[27] = 1'b1;
      zz_rom_89[28] = 1'b1;
      zz_rom_89[29] = 1'b1;
      zz_rom_89[30] = 1'b1;
      zz_rom_89[31] = 1'b1;
      zz_rom_89[32] = 1'b1;
      zz_rom_89[33] = 1'b1;
      zz_rom_89[34] = 1'b1;
      zz_rom_89[35] = 1'b1;
      zz_rom_89[36] = 1'b1;
      zz_rom_89[37] = 1'b1;
      zz_rom_89[38] = 1'b1;
      zz_rom_89[39] = 1'b1;
      zz_rom_89[40] = 1'b1;
      zz_rom_89[41] = 1'b1;
      zz_rom_89[42] = 1'b1;
      zz_rom_89[43] = 1'b1;
      zz_rom_89[44] = 1'b1;
      zz_rom_89[45] = 1'b1;
      zz_rom_89[46] = 1'b1;
      zz_rom_89[47] = 1'b1;
      zz_rom_89[48] = 1'b1;
      zz_rom_89[49] = 1'b1;
      zz_rom_89[50] = 1'b1;
      zz_rom_89[51] = 1'b1;
      zz_rom_89[52] = 1'b1;
      zz_rom_89[53] = 1'b1;
      zz_rom_89[54] = 1'b1;
      zz_rom_89[55] = 1'b1;
      zz_rom_89[56] = 1'b1;
      zz_rom_89[57] = 1'b1;
      zz_rom_89[58] = 1'b1;
      zz_rom_89[59] = 1'b1;
      zz_rom_89[60] = 1'b1;
      zz_rom_89[61] = 1'b1;
      zz_rom_89[62] = 1'b1;
      zz_rom_89[63] = 1'b1;
      zz_rom_89[64] = 1'b1;
      zz_rom_89[65] = 1'b1;
      zz_rom_89[66] = 1'b1;
      zz_rom_89[67] = 1'b1;
      zz_rom_89[68] = 1'b1;
      zz_rom_89[69] = 1'b1;
      zz_rom_89[70] = 1'b1;
      zz_rom_89[71] = 1'b1;
      zz_rom_89[72] = 1'b1;
      zz_rom_89[73] = 1'b1;
      zz_rom_89[74] = 1'b1;
      zz_rom_89[75] = 1'b1;
      zz_rom_89[76] = 1'b1;
      zz_rom_89[77] = 1'b1;
      zz_rom_89[78] = 1'b1;
      zz_rom_89[79] = 1'b1;
      zz_rom_89[80] = 1'b1;
      zz_rom_89[81] = 1'b1;
      zz_rom_89[82] = 1'b0;
      zz_rom_89[83] = 1'b0;
      zz_rom_89[84] = 1'b0;
      zz_rom_89[85] = 1'b0;
      zz_rom_89[86] = 1'b0;
      zz_rom_89[87] = 1'b0;
      zz_rom_89[88] = 1'b0;
      zz_rom_89[89] = 1'b0;
      zz_rom_89[90] = 1'b0;
      zz_rom_89[91] = 1'b0;
      zz_rom_89[92] = 1'b0;
      zz_rom_89[93] = 1'b0;
      zz_rom_89[94] = 1'b0;
      zz_rom_89[95] = 1'b0;
      zz_rom_89[96] = 1'b0;
      zz_rom_89[97] = 1'b0;
      zz_rom_89[98] = 1'b0;
      zz_rom_89[99] = 1'b0;
    end
  endfunction
  wire [99:0] _zz_90;
  function [99:0] zz_rom_90(input dummy);
    begin
      zz_rom_90[0] = 1'b0;
      zz_rom_90[1] = 1'b0;
      zz_rom_90[2] = 1'b0;
      zz_rom_90[3] = 1'b0;
      zz_rom_90[4] = 1'b0;
      zz_rom_90[5] = 1'b0;
      zz_rom_90[6] = 1'b0;
      zz_rom_90[7] = 1'b0;
      zz_rom_90[8] = 1'b0;
      zz_rom_90[9] = 1'b0;
      zz_rom_90[10] = 1'b0;
      zz_rom_90[11] = 1'b0;
      zz_rom_90[12] = 1'b0;
      zz_rom_90[13] = 1'b0;
      zz_rom_90[14] = 1'b0;
      zz_rom_90[15] = 1'b0;
      zz_rom_90[16] = 1'b0;
      zz_rom_90[17] = 1'b0;
      zz_rom_90[18] = 1'b0;
      zz_rom_90[19] = 1'b0;
      zz_rom_90[20] = 1'b1;
      zz_rom_90[21] = 1'b1;
      zz_rom_90[22] = 1'b1;
      zz_rom_90[23] = 1'b1;
      zz_rom_90[24] = 1'b1;
      zz_rom_90[25] = 1'b1;
      zz_rom_90[26] = 1'b1;
      zz_rom_90[27] = 1'b1;
      zz_rom_90[28] = 1'b1;
      zz_rom_90[29] = 1'b1;
      zz_rom_90[30] = 1'b1;
      zz_rom_90[31] = 1'b1;
      zz_rom_90[32] = 1'b1;
      zz_rom_90[33] = 1'b1;
      zz_rom_90[34] = 1'b1;
      zz_rom_90[35] = 1'b1;
      zz_rom_90[36] = 1'b1;
      zz_rom_90[37] = 1'b1;
      zz_rom_90[38] = 1'b1;
      zz_rom_90[39] = 1'b1;
      zz_rom_90[40] = 1'b1;
      zz_rom_90[41] = 1'b1;
      zz_rom_90[42] = 1'b1;
      zz_rom_90[43] = 1'b1;
      zz_rom_90[44] = 1'b1;
      zz_rom_90[45] = 1'b1;
      zz_rom_90[46] = 1'b1;
      zz_rom_90[47] = 1'b1;
      zz_rom_90[48] = 1'b1;
      zz_rom_90[49] = 1'b1;
      zz_rom_90[50] = 1'b1;
      zz_rom_90[51] = 1'b1;
      zz_rom_90[52] = 1'b1;
      zz_rom_90[53] = 1'b1;
      zz_rom_90[54] = 1'b1;
      zz_rom_90[55] = 1'b1;
      zz_rom_90[56] = 1'b1;
      zz_rom_90[57] = 1'b1;
      zz_rom_90[58] = 1'b1;
      zz_rom_90[59] = 1'b1;
      zz_rom_90[60] = 1'b1;
      zz_rom_90[61] = 1'b1;
      zz_rom_90[62] = 1'b1;
      zz_rom_90[63] = 1'b1;
      zz_rom_90[64] = 1'b1;
      zz_rom_90[65] = 1'b1;
      zz_rom_90[66] = 1'b1;
      zz_rom_90[67] = 1'b1;
      zz_rom_90[68] = 1'b1;
      zz_rom_90[69] = 1'b1;
      zz_rom_90[70] = 1'b1;
      zz_rom_90[71] = 1'b1;
      zz_rom_90[72] = 1'b1;
      zz_rom_90[73] = 1'b1;
      zz_rom_90[74] = 1'b1;
      zz_rom_90[75] = 1'b1;
      zz_rom_90[76] = 1'b1;
      zz_rom_90[77] = 1'b1;
      zz_rom_90[78] = 1'b1;
      zz_rom_90[79] = 1'b1;
      zz_rom_90[80] = 1'b1;
      zz_rom_90[81] = 1'b0;
      zz_rom_90[82] = 1'b0;
      zz_rom_90[83] = 1'b0;
      zz_rom_90[84] = 1'b0;
      zz_rom_90[85] = 1'b0;
      zz_rom_90[86] = 1'b0;
      zz_rom_90[87] = 1'b0;
      zz_rom_90[88] = 1'b0;
      zz_rom_90[89] = 1'b0;
      zz_rom_90[90] = 1'b0;
      zz_rom_90[91] = 1'b0;
      zz_rom_90[92] = 1'b0;
      zz_rom_90[93] = 1'b0;
      zz_rom_90[94] = 1'b0;
      zz_rom_90[95] = 1'b0;
      zz_rom_90[96] = 1'b0;
      zz_rom_90[97] = 1'b0;
      zz_rom_90[98] = 1'b0;
      zz_rom_90[99] = 1'b0;
    end
  endfunction
  wire [99:0] _zz_91;
  function [99:0] zz_rom_91(input dummy);
    begin
      zz_rom_91[0] = 1'b0;
      zz_rom_91[1] = 1'b0;
      zz_rom_91[2] = 1'b0;
      zz_rom_91[3] = 1'b0;
      zz_rom_91[4] = 1'b0;
      zz_rom_91[5] = 1'b0;
      zz_rom_91[6] = 1'b0;
      zz_rom_91[7] = 1'b0;
      zz_rom_91[8] = 1'b0;
      zz_rom_91[9] = 1'b0;
      zz_rom_91[10] = 1'b0;
      zz_rom_91[11] = 1'b0;
      zz_rom_91[12] = 1'b0;
      zz_rom_91[13] = 1'b0;
      zz_rom_91[14] = 1'b0;
      zz_rom_91[15] = 1'b0;
      zz_rom_91[16] = 1'b0;
      zz_rom_91[17] = 1'b0;
      zz_rom_91[18] = 1'b0;
      zz_rom_91[19] = 1'b0;
      zz_rom_91[20] = 1'b0;
      zz_rom_91[21] = 1'b0;
      zz_rom_91[22] = 1'b1;
      zz_rom_91[23] = 1'b1;
      zz_rom_91[24] = 1'b1;
      zz_rom_91[25] = 1'b1;
      zz_rom_91[26] = 1'b1;
      zz_rom_91[27] = 1'b1;
      zz_rom_91[28] = 1'b1;
      zz_rom_91[29] = 1'b1;
      zz_rom_91[30] = 1'b1;
      zz_rom_91[31] = 1'b1;
      zz_rom_91[32] = 1'b1;
      zz_rom_91[33] = 1'b1;
      zz_rom_91[34] = 1'b1;
      zz_rom_91[35] = 1'b1;
      zz_rom_91[36] = 1'b1;
      zz_rom_91[37] = 1'b1;
      zz_rom_91[38] = 1'b1;
      zz_rom_91[39] = 1'b1;
      zz_rom_91[40] = 1'b1;
      zz_rom_91[41] = 1'b1;
      zz_rom_91[42] = 1'b1;
      zz_rom_91[43] = 1'b1;
      zz_rom_91[44] = 1'b1;
      zz_rom_91[45] = 1'b1;
      zz_rom_91[46] = 1'b1;
      zz_rom_91[47] = 1'b1;
      zz_rom_91[48] = 1'b1;
      zz_rom_91[49] = 1'b1;
      zz_rom_91[50] = 1'b1;
      zz_rom_91[51] = 1'b1;
      zz_rom_91[52] = 1'b1;
      zz_rom_91[53] = 1'b1;
      zz_rom_91[54] = 1'b1;
      zz_rom_91[55] = 1'b1;
      zz_rom_91[56] = 1'b1;
      zz_rom_91[57] = 1'b1;
      zz_rom_91[58] = 1'b1;
      zz_rom_91[59] = 1'b1;
      zz_rom_91[60] = 1'b1;
      zz_rom_91[61] = 1'b1;
      zz_rom_91[62] = 1'b1;
      zz_rom_91[63] = 1'b1;
      zz_rom_91[64] = 1'b1;
      zz_rom_91[65] = 1'b1;
      zz_rom_91[66] = 1'b1;
      zz_rom_91[67] = 1'b1;
      zz_rom_91[68] = 1'b1;
      zz_rom_91[69] = 1'b1;
      zz_rom_91[70] = 1'b1;
      zz_rom_91[71] = 1'b1;
      zz_rom_91[72] = 1'b1;
      zz_rom_91[73] = 1'b1;
      zz_rom_91[74] = 1'b1;
      zz_rom_91[75] = 1'b1;
      zz_rom_91[76] = 1'b1;
      zz_rom_91[77] = 1'b1;
      zz_rom_91[78] = 1'b1;
      zz_rom_91[79] = 1'b0;
      zz_rom_91[80] = 1'b0;
      zz_rom_91[81] = 1'b0;
      zz_rom_91[82] = 1'b0;
      zz_rom_91[83] = 1'b0;
      zz_rom_91[84] = 1'b0;
      zz_rom_91[85] = 1'b0;
      zz_rom_91[86] = 1'b0;
      zz_rom_91[87] = 1'b0;
      zz_rom_91[88] = 1'b0;
      zz_rom_91[89] = 1'b0;
      zz_rom_91[90] = 1'b0;
      zz_rom_91[91] = 1'b0;
      zz_rom_91[92] = 1'b0;
      zz_rom_91[93] = 1'b0;
      zz_rom_91[94] = 1'b0;
      zz_rom_91[95] = 1'b0;
      zz_rom_91[96] = 1'b0;
      zz_rom_91[97] = 1'b0;
      zz_rom_91[98] = 1'b0;
      zz_rom_91[99] = 1'b0;
    end
  endfunction
  wire [99:0] _zz_92;
  function [99:0] zz_rom_92(input dummy);
    begin
      zz_rom_92[0] = 1'b0;
      zz_rom_92[1] = 1'b0;
      zz_rom_92[2] = 1'b0;
      zz_rom_92[3] = 1'b0;
      zz_rom_92[4] = 1'b0;
      zz_rom_92[5] = 1'b0;
      zz_rom_92[6] = 1'b0;
      zz_rom_92[7] = 1'b0;
      zz_rom_92[8] = 1'b0;
      zz_rom_92[9] = 1'b0;
      zz_rom_92[10] = 1'b0;
      zz_rom_92[11] = 1'b0;
      zz_rom_92[12] = 1'b0;
      zz_rom_92[13] = 1'b0;
      zz_rom_92[14] = 1'b0;
      zz_rom_92[15] = 1'b0;
      zz_rom_92[16] = 1'b0;
      zz_rom_92[17] = 1'b0;
      zz_rom_92[18] = 1'b0;
      zz_rom_92[19] = 1'b0;
      zz_rom_92[20] = 1'b0;
      zz_rom_92[21] = 1'b0;
      zz_rom_92[22] = 1'b0;
      zz_rom_92[23] = 1'b1;
      zz_rom_92[24] = 1'b1;
      zz_rom_92[25] = 1'b1;
      zz_rom_92[26] = 1'b1;
      zz_rom_92[27] = 1'b1;
      zz_rom_92[28] = 1'b1;
      zz_rom_92[29] = 1'b1;
      zz_rom_92[30] = 1'b1;
      zz_rom_92[31] = 1'b1;
      zz_rom_92[32] = 1'b1;
      zz_rom_92[33] = 1'b1;
      zz_rom_92[34] = 1'b1;
      zz_rom_92[35] = 1'b1;
      zz_rom_92[36] = 1'b1;
      zz_rom_92[37] = 1'b1;
      zz_rom_92[38] = 1'b1;
      zz_rom_92[39] = 1'b1;
      zz_rom_92[40] = 1'b1;
      zz_rom_92[41] = 1'b1;
      zz_rom_92[42] = 1'b1;
      zz_rom_92[43] = 1'b1;
      zz_rom_92[44] = 1'b1;
      zz_rom_92[45] = 1'b1;
      zz_rom_92[46] = 1'b1;
      zz_rom_92[47] = 1'b1;
      zz_rom_92[48] = 1'b1;
      zz_rom_92[49] = 1'b1;
      zz_rom_92[50] = 1'b1;
      zz_rom_92[51] = 1'b1;
      zz_rom_92[52] = 1'b1;
      zz_rom_92[53] = 1'b1;
      zz_rom_92[54] = 1'b1;
      zz_rom_92[55] = 1'b1;
      zz_rom_92[56] = 1'b1;
      zz_rom_92[57] = 1'b1;
      zz_rom_92[58] = 1'b1;
      zz_rom_92[59] = 1'b1;
      zz_rom_92[60] = 1'b1;
      zz_rom_92[61] = 1'b1;
      zz_rom_92[62] = 1'b1;
      zz_rom_92[63] = 1'b1;
      zz_rom_92[64] = 1'b1;
      zz_rom_92[65] = 1'b1;
      zz_rom_92[66] = 1'b1;
      zz_rom_92[67] = 1'b1;
      zz_rom_92[68] = 1'b1;
      zz_rom_92[69] = 1'b1;
      zz_rom_92[70] = 1'b1;
      zz_rom_92[71] = 1'b1;
      zz_rom_92[72] = 1'b1;
      zz_rom_92[73] = 1'b1;
      zz_rom_92[74] = 1'b1;
      zz_rom_92[75] = 1'b1;
      zz_rom_92[76] = 1'b1;
      zz_rom_92[77] = 1'b1;
      zz_rom_92[78] = 1'b0;
      zz_rom_92[79] = 1'b0;
      zz_rom_92[80] = 1'b0;
      zz_rom_92[81] = 1'b0;
      zz_rom_92[82] = 1'b0;
      zz_rom_92[83] = 1'b0;
      zz_rom_92[84] = 1'b0;
      zz_rom_92[85] = 1'b0;
      zz_rom_92[86] = 1'b0;
      zz_rom_92[87] = 1'b0;
      zz_rom_92[88] = 1'b0;
      zz_rom_92[89] = 1'b0;
      zz_rom_92[90] = 1'b0;
      zz_rom_92[91] = 1'b0;
      zz_rom_92[92] = 1'b0;
      zz_rom_92[93] = 1'b0;
      zz_rom_92[94] = 1'b0;
      zz_rom_92[95] = 1'b0;
      zz_rom_92[96] = 1'b0;
      zz_rom_92[97] = 1'b0;
      zz_rom_92[98] = 1'b0;
      zz_rom_92[99] = 1'b0;
    end
  endfunction
  wire [99:0] _zz_93;
  function [99:0] zz_rom_93(input dummy);
    begin
      zz_rom_93[0] = 1'b0;
      zz_rom_93[1] = 1'b0;
      zz_rom_93[2] = 1'b0;
      zz_rom_93[3] = 1'b0;
      zz_rom_93[4] = 1'b0;
      zz_rom_93[5] = 1'b0;
      zz_rom_93[6] = 1'b0;
      zz_rom_93[7] = 1'b0;
      zz_rom_93[8] = 1'b0;
      zz_rom_93[9] = 1'b0;
      zz_rom_93[10] = 1'b0;
      zz_rom_93[11] = 1'b0;
      zz_rom_93[12] = 1'b0;
      zz_rom_93[13] = 1'b0;
      zz_rom_93[14] = 1'b0;
      zz_rom_93[15] = 1'b0;
      zz_rom_93[16] = 1'b0;
      zz_rom_93[17] = 1'b0;
      zz_rom_93[18] = 1'b0;
      zz_rom_93[19] = 1'b0;
      zz_rom_93[20] = 1'b0;
      zz_rom_93[21] = 1'b0;
      zz_rom_93[22] = 1'b0;
      zz_rom_93[23] = 1'b0;
      zz_rom_93[24] = 1'b0;
      zz_rom_93[25] = 1'b1;
      zz_rom_93[26] = 1'b1;
      zz_rom_93[27] = 1'b1;
      zz_rom_93[28] = 1'b1;
      zz_rom_93[29] = 1'b1;
      zz_rom_93[30] = 1'b1;
      zz_rom_93[31] = 1'b1;
      zz_rom_93[32] = 1'b1;
      zz_rom_93[33] = 1'b1;
      zz_rom_93[34] = 1'b1;
      zz_rom_93[35] = 1'b1;
      zz_rom_93[36] = 1'b1;
      zz_rom_93[37] = 1'b1;
      zz_rom_93[38] = 1'b1;
      zz_rom_93[39] = 1'b1;
      zz_rom_93[40] = 1'b1;
      zz_rom_93[41] = 1'b1;
      zz_rom_93[42] = 1'b1;
      zz_rom_93[43] = 1'b1;
      zz_rom_93[44] = 1'b1;
      zz_rom_93[45] = 1'b1;
      zz_rom_93[46] = 1'b1;
      zz_rom_93[47] = 1'b1;
      zz_rom_93[48] = 1'b1;
      zz_rom_93[49] = 1'b1;
      zz_rom_93[50] = 1'b1;
      zz_rom_93[51] = 1'b1;
      zz_rom_93[52] = 1'b1;
      zz_rom_93[53] = 1'b1;
      zz_rom_93[54] = 1'b1;
      zz_rom_93[55] = 1'b1;
      zz_rom_93[56] = 1'b1;
      zz_rom_93[57] = 1'b1;
      zz_rom_93[58] = 1'b1;
      zz_rom_93[59] = 1'b1;
      zz_rom_93[60] = 1'b1;
      zz_rom_93[61] = 1'b1;
      zz_rom_93[62] = 1'b1;
      zz_rom_93[63] = 1'b1;
      zz_rom_93[64] = 1'b1;
      zz_rom_93[65] = 1'b1;
      zz_rom_93[66] = 1'b1;
      zz_rom_93[67] = 1'b1;
      zz_rom_93[68] = 1'b1;
      zz_rom_93[69] = 1'b1;
      zz_rom_93[70] = 1'b1;
      zz_rom_93[71] = 1'b1;
      zz_rom_93[72] = 1'b1;
      zz_rom_93[73] = 1'b1;
      zz_rom_93[74] = 1'b1;
      zz_rom_93[75] = 1'b1;
      zz_rom_93[76] = 1'b0;
      zz_rom_93[77] = 1'b0;
      zz_rom_93[78] = 1'b0;
      zz_rom_93[79] = 1'b0;
      zz_rom_93[80] = 1'b0;
      zz_rom_93[81] = 1'b0;
      zz_rom_93[82] = 1'b0;
      zz_rom_93[83] = 1'b0;
      zz_rom_93[84] = 1'b0;
      zz_rom_93[85] = 1'b0;
      zz_rom_93[86] = 1'b0;
      zz_rom_93[87] = 1'b0;
      zz_rom_93[88] = 1'b0;
      zz_rom_93[89] = 1'b0;
      zz_rom_93[90] = 1'b0;
      zz_rom_93[91] = 1'b0;
      zz_rom_93[92] = 1'b0;
      zz_rom_93[93] = 1'b0;
      zz_rom_93[94] = 1'b0;
      zz_rom_93[95] = 1'b0;
      zz_rom_93[96] = 1'b0;
      zz_rom_93[97] = 1'b0;
      zz_rom_93[98] = 1'b0;
      zz_rom_93[99] = 1'b0;
    end
  endfunction
  wire [99:0] _zz_94;
  function [99:0] zz_rom_94(input dummy);
    begin
      zz_rom_94[0] = 1'b0;
      zz_rom_94[1] = 1'b0;
      zz_rom_94[2] = 1'b0;
      zz_rom_94[3] = 1'b0;
      zz_rom_94[4] = 1'b0;
      zz_rom_94[5] = 1'b0;
      zz_rom_94[6] = 1'b0;
      zz_rom_94[7] = 1'b0;
      zz_rom_94[8] = 1'b0;
      zz_rom_94[9] = 1'b0;
      zz_rom_94[10] = 1'b0;
      zz_rom_94[11] = 1'b0;
      zz_rom_94[12] = 1'b0;
      zz_rom_94[13] = 1'b0;
      zz_rom_94[14] = 1'b0;
      zz_rom_94[15] = 1'b0;
      zz_rom_94[16] = 1'b0;
      zz_rom_94[17] = 1'b0;
      zz_rom_94[18] = 1'b0;
      zz_rom_94[19] = 1'b0;
      zz_rom_94[20] = 1'b0;
      zz_rom_94[21] = 1'b0;
      zz_rom_94[22] = 1'b0;
      zz_rom_94[23] = 1'b0;
      zz_rom_94[24] = 1'b0;
      zz_rom_94[25] = 1'b0;
      zz_rom_94[26] = 1'b0;
      zz_rom_94[27] = 1'b1;
      zz_rom_94[28] = 1'b1;
      zz_rom_94[29] = 1'b1;
      zz_rom_94[30] = 1'b1;
      zz_rom_94[31] = 1'b1;
      zz_rom_94[32] = 1'b1;
      zz_rom_94[33] = 1'b1;
      zz_rom_94[34] = 1'b1;
      zz_rom_94[35] = 1'b1;
      zz_rom_94[36] = 1'b1;
      zz_rom_94[37] = 1'b1;
      zz_rom_94[38] = 1'b1;
      zz_rom_94[39] = 1'b1;
      zz_rom_94[40] = 1'b1;
      zz_rom_94[41] = 1'b1;
      zz_rom_94[42] = 1'b1;
      zz_rom_94[43] = 1'b1;
      zz_rom_94[44] = 1'b1;
      zz_rom_94[45] = 1'b1;
      zz_rom_94[46] = 1'b1;
      zz_rom_94[47] = 1'b1;
      zz_rom_94[48] = 1'b1;
      zz_rom_94[49] = 1'b1;
      zz_rom_94[50] = 1'b1;
      zz_rom_94[51] = 1'b1;
      zz_rom_94[52] = 1'b1;
      zz_rom_94[53] = 1'b1;
      zz_rom_94[54] = 1'b1;
      zz_rom_94[55] = 1'b1;
      zz_rom_94[56] = 1'b1;
      zz_rom_94[57] = 1'b1;
      zz_rom_94[58] = 1'b1;
      zz_rom_94[59] = 1'b1;
      zz_rom_94[60] = 1'b1;
      zz_rom_94[61] = 1'b1;
      zz_rom_94[62] = 1'b1;
      zz_rom_94[63] = 1'b1;
      zz_rom_94[64] = 1'b1;
      zz_rom_94[65] = 1'b1;
      zz_rom_94[66] = 1'b1;
      zz_rom_94[67] = 1'b1;
      zz_rom_94[68] = 1'b1;
      zz_rom_94[69] = 1'b1;
      zz_rom_94[70] = 1'b1;
      zz_rom_94[71] = 1'b1;
      zz_rom_94[72] = 1'b1;
      zz_rom_94[73] = 1'b1;
      zz_rom_94[74] = 1'b0;
      zz_rom_94[75] = 1'b0;
      zz_rom_94[76] = 1'b0;
      zz_rom_94[77] = 1'b0;
      zz_rom_94[78] = 1'b0;
      zz_rom_94[79] = 1'b0;
      zz_rom_94[80] = 1'b0;
      zz_rom_94[81] = 1'b0;
      zz_rom_94[82] = 1'b0;
      zz_rom_94[83] = 1'b0;
      zz_rom_94[84] = 1'b0;
      zz_rom_94[85] = 1'b0;
      zz_rom_94[86] = 1'b0;
      zz_rom_94[87] = 1'b0;
      zz_rom_94[88] = 1'b0;
      zz_rom_94[89] = 1'b0;
      zz_rom_94[90] = 1'b0;
      zz_rom_94[91] = 1'b0;
      zz_rom_94[92] = 1'b0;
      zz_rom_94[93] = 1'b0;
      zz_rom_94[94] = 1'b0;
      zz_rom_94[95] = 1'b0;
      zz_rom_94[96] = 1'b0;
      zz_rom_94[97] = 1'b0;
      zz_rom_94[98] = 1'b0;
      zz_rom_94[99] = 1'b0;
    end
  endfunction
  wire [99:0] _zz_95;
  function [99:0] zz_rom_95(input dummy);
    begin
      zz_rom_95[0] = 1'b0;
      zz_rom_95[1] = 1'b0;
      zz_rom_95[2] = 1'b0;
      zz_rom_95[3] = 1'b0;
      zz_rom_95[4] = 1'b0;
      zz_rom_95[5] = 1'b0;
      zz_rom_95[6] = 1'b0;
      zz_rom_95[7] = 1'b0;
      zz_rom_95[8] = 1'b0;
      zz_rom_95[9] = 1'b0;
      zz_rom_95[10] = 1'b0;
      zz_rom_95[11] = 1'b0;
      zz_rom_95[12] = 1'b0;
      zz_rom_95[13] = 1'b0;
      zz_rom_95[14] = 1'b0;
      zz_rom_95[15] = 1'b0;
      zz_rom_95[16] = 1'b0;
      zz_rom_95[17] = 1'b0;
      zz_rom_95[18] = 1'b0;
      zz_rom_95[19] = 1'b0;
      zz_rom_95[20] = 1'b0;
      zz_rom_95[21] = 1'b0;
      zz_rom_95[22] = 1'b0;
      zz_rom_95[23] = 1'b0;
      zz_rom_95[24] = 1'b0;
      zz_rom_95[25] = 1'b0;
      zz_rom_95[26] = 1'b0;
      zz_rom_95[27] = 1'b0;
      zz_rom_95[28] = 1'b0;
      zz_rom_95[29] = 1'b1;
      zz_rom_95[30] = 1'b1;
      zz_rom_95[31] = 1'b1;
      zz_rom_95[32] = 1'b1;
      zz_rom_95[33] = 1'b1;
      zz_rom_95[34] = 1'b1;
      zz_rom_95[35] = 1'b1;
      zz_rom_95[36] = 1'b1;
      zz_rom_95[37] = 1'b1;
      zz_rom_95[38] = 1'b1;
      zz_rom_95[39] = 1'b1;
      zz_rom_95[40] = 1'b1;
      zz_rom_95[41] = 1'b1;
      zz_rom_95[42] = 1'b1;
      zz_rom_95[43] = 1'b1;
      zz_rom_95[44] = 1'b1;
      zz_rom_95[45] = 1'b1;
      zz_rom_95[46] = 1'b1;
      zz_rom_95[47] = 1'b1;
      zz_rom_95[48] = 1'b1;
      zz_rom_95[49] = 1'b1;
      zz_rom_95[50] = 1'b1;
      zz_rom_95[51] = 1'b1;
      zz_rom_95[52] = 1'b1;
      zz_rom_95[53] = 1'b1;
      zz_rom_95[54] = 1'b1;
      zz_rom_95[55] = 1'b1;
      zz_rom_95[56] = 1'b1;
      zz_rom_95[57] = 1'b1;
      zz_rom_95[58] = 1'b1;
      zz_rom_95[59] = 1'b1;
      zz_rom_95[60] = 1'b1;
      zz_rom_95[61] = 1'b1;
      zz_rom_95[62] = 1'b1;
      zz_rom_95[63] = 1'b1;
      zz_rom_95[64] = 1'b1;
      zz_rom_95[65] = 1'b1;
      zz_rom_95[66] = 1'b1;
      zz_rom_95[67] = 1'b1;
      zz_rom_95[68] = 1'b1;
      zz_rom_95[69] = 1'b1;
      zz_rom_95[70] = 1'b1;
      zz_rom_95[71] = 1'b1;
      zz_rom_95[72] = 1'b0;
      zz_rom_95[73] = 1'b0;
      zz_rom_95[74] = 1'b0;
      zz_rom_95[75] = 1'b0;
      zz_rom_95[76] = 1'b0;
      zz_rom_95[77] = 1'b0;
      zz_rom_95[78] = 1'b0;
      zz_rom_95[79] = 1'b0;
      zz_rom_95[80] = 1'b0;
      zz_rom_95[81] = 1'b0;
      zz_rom_95[82] = 1'b0;
      zz_rom_95[83] = 1'b0;
      zz_rom_95[84] = 1'b0;
      zz_rom_95[85] = 1'b0;
      zz_rom_95[86] = 1'b0;
      zz_rom_95[87] = 1'b0;
      zz_rom_95[88] = 1'b0;
      zz_rom_95[89] = 1'b0;
      zz_rom_95[90] = 1'b0;
      zz_rom_95[91] = 1'b0;
      zz_rom_95[92] = 1'b0;
      zz_rom_95[93] = 1'b0;
      zz_rom_95[94] = 1'b0;
      zz_rom_95[95] = 1'b0;
      zz_rom_95[96] = 1'b0;
      zz_rom_95[97] = 1'b0;
      zz_rom_95[98] = 1'b0;
      zz_rom_95[99] = 1'b0;
    end
  endfunction
  wire [99:0] _zz_96;
  function [99:0] zz_rom_96(input dummy);
    begin
      zz_rom_96[0] = 1'b0;
      zz_rom_96[1] = 1'b0;
      zz_rom_96[2] = 1'b0;
      zz_rom_96[3] = 1'b0;
      zz_rom_96[4] = 1'b0;
      zz_rom_96[5] = 1'b0;
      zz_rom_96[6] = 1'b0;
      zz_rom_96[7] = 1'b0;
      zz_rom_96[8] = 1'b0;
      zz_rom_96[9] = 1'b0;
      zz_rom_96[10] = 1'b0;
      zz_rom_96[11] = 1'b0;
      zz_rom_96[12] = 1'b0;
      zz_rom_96[13] = 1'b0;
      zz_rom_96[14] = 1'b0;
      zz_rom_96[15] = 1'b0;
      zz_rom_96[16] = 1'b0;
      zz_rom_96[17] = 1'b0;
      zz_rom_96[18] = 1'b0;
      zz_rom_96[19] = 1'b0;
      zz_rom_96[20] = 1'b0;
      zz_rom_96[21] = 1'b0;
      zz_rom_96[22] = 1'b0;
      zz_rom_96[23] = 1'b0;
      zz_rom_96[24] = 1'b0;
      zz_rom_96[25] = 1'b0;
      zz_rom_96[26] = 1'b0;
      zz_rom_96[27] = 1'b0;
      zz_rom_96[28] = 1'b0;
      zz_rom_96[29] = 1'b0;
      zz_rom_96[30] = 1'b0;
      zz_rom_96[31] = 1'b1;
      zz_rom_96[32] = 1'b1;
      zz_rom_96[33] = 1'b1;
      zz_rom_96[34] = 1'b1;
      zz_rom_96[35] = 1'b1;
      zz_rom_96[36] = 1'b1;
      zz_rom_96[37] = 1'b1;
      zz_rom_96[38] = 1'b1;
      zz_rom_96[39] = 1'b1;
      zz_rom_96[40] = 1'b1;
      zz_rom_96[41] = 1'b1;
      zz_rom_96[42] = 1'b1;
      zz_rom_96[43] = 1'b1;
      zz_rom_96[44] = 1'b1;
      zz_rom_96[45] = 1'b1;
      zz_rom_96[46] = 1'b1;
      zz_rom_96[47] = 1'b1;
      zz_rom_96[48] = 1'b1;
      zz_rom_96[49] = 1'b1;
      zz_rom_96[50] = 1'b1;
      zz_rom_96[51] = 1'b1;
      zz_rom_96[52] = 1'b1;
      zz_rom_96[53] = 1'b1;
      zz_rom_96[54] = 1'b1;
      zz_rom_96[55] = 1'b1;
      zz_rom_96[56] = 1'b1;
      zz_rom_96[57] = 1'b1;
      zz_rom_96[58] = 1'b1;
      zz_rom_96[59] = 1'b1;
      zz_rom_96[60] = 1'b1;
      zz_rom_96[61] = 1'b1;
      zz_rom_96[62] = 1'b1;
      zz_rom_96[63] = 1'b1;
      zz_rom_96[64] = 1'b1;
      zz_rom_96[65] = 1'b1;
      zz_rom_96[66] = 1'b1;
      zz_rom_96[67] = 1'b1;
      zz_rom_96[68] = 1'b1;
      zz_rom_96[69] = 1'b1;
      zz_rom_96[70] = 1'b0;
      zz_rom_96[71] = 1'b0;
      zz_rom_96[72] = 1'b0;
      zz_rom_96[73] = 1'b0;
      zz_rom_96[74] = 1'b0;
      zz_rom_96[75] = 1'b0;
      zz_rom_96[76] = 1'b0;
      zz_rom_96[77] = 1'b0;
      zz_rom_96[78] = 1'b0;
      zz_rom_96[79] = 1'b0;
      zz_rom_96[80] = 1'b0;
      zz_rom_96[81] = 1'b0;
      zz_rom_96[82] = 1'b0;
      zz_rom_96[83] = 1'b0;
      zz_rom_96[84] = 1'b0;
      zz_rom_96[85] = 1'b0;
      zz_rom_96[86] = 1'b0;
      zz_rom_96[87] = 1'b0;
      zz_rom_96[88] = 1'b0;
      zz_rom_96[89] = 1'b0;
      zz_rom_96[90] = 1'b0;
      zz_rom_96[91] = 1'b0;
      zz_rom_96[92] = 1'b0;
      zz_rom_96[93] = 1'b0;
      zz_rom_96[94] = 1'b0;
      zz_rom_96[95] = 1'b0;
      zz_rom_96[96] = 1'b0;
      zz_rom_96[97] = 1'b0;
      zz_rom_96[98] = 1'b0;
      zz_rom_96[99] = 1'b0;
    end
  endfunction
  wire [99:0] _zz_97;
  function [99:0] zz_rom_97(input dummy);
    begin
      zz_rom_97[0] = 1'b0;
      zz_rom_97[1] = 1'b0;
      zz_rom_97[2] = 1'b0;
      zz_rom_97[3] = 1'b0;
      zz_rom_97[4] = 1'b0;
      zz_rom_97[5] = 1'b0;
      zz_rom_97[6] = 1'b0;
      zz_rom_97[7] = 1'b0;
      zz_rom_97[8] = 1'b0;
      zz_rom_97[9] = 1'b0;
      zz_rom_97[10] = 1'b0;
      zz_rom_97[11] = 1'b0;
      zz_rom_97[12] = 1'b0;
      zz_rom_97[13] = 1'b0;
      zz_rom_97[14] = 1'b0;
      zz_rom_97[15] = 1'b0;
      zz_rom_97[16] = 1'b0;
      zz_rom_97[17] = 1'b0;
      zz_rom_97[18] = 1'b0;
      zz_rom_97[19] = 1'b0;
      zz_rom_97[20] = 1'b0;
      zz_rom_97[21] = 1'b0;
      zz_rom_97[22] = 1'b0;
      zz_rom_97[23] = 1'b0;
      zz_rom_97[24] = 1'b0;
      zz_rom_97[25] = 1'b0;
      zz_rom_97[26] = 1'b0;
      zz_rom_97[27] = 1'b0;
      zz_rom_97[28] = 1'b0;
      zz_rom_97[29] = 1'b0;
      zz_rom_97[30] = 1'b0;
      zz_rom_97[31] = 1'b0;
      zz_rom_97[32] = 1'b0;
      zz_rom_97[33] = 1'b1;
      zz_rom_97[34] = 1'b1;
      zz_rom_97[35] = 1'b1;
      zz_rom_97[36] = 1'b1;
      zz_rom_97[37] = 1'b1;
      zz_rom_97[38] = 1'b1;
      zz_rom_97[39] = 1'b1;
      zz_rom_97[40] = 1'b1;
      zz_rom_97[41] = 1'b1;
      zz_rom_97[42] = 1'b1;
      zz_rom_97[43] = 1'b1;
      zz_rom_97[44] = 1'b1;
      zz_rom_97[45] = 1'b1;
      zz_rom_97[46] = 1'b1;
      zz_rom_97[47] = 1'b1;
      zz_rom_97[48] = 1'b1;
      zz_rom_97[49] = 1'b1;
      zz_rom_97[50] = 1'b1;
      zz_rom_97[51] = 1'b1;
      zz_rom_97[52] = 1'b1;
      zz_rom_97[53] = 1'b1;
      zz_rom_97[54] = 1'b1;
      zz_rom_97[55] = 1'b1;
      zz_rom_97[56] = 1'b1;
      zz_rom_97[57] = 1'b1;
      zz_rom_97[58] = 1'b1;
      zz_rom_97[59] = 1'b1;
      zz_rom_97[60] = 1'b1;
      zz_rom_97[61] = 1'b1;
      zz_rom_97[62] = 1'b1;
      zz_rom_97[63] = 1'b1;
      zz_rom_97[64] = 1'b1;
      zz_rom_97[65] = 1'b1;
      zz_rom_97[66] = 1'b1;
      zz_rom_97[67] = 1'b1;
      zz_rom_97[68] = 1'b0;
      zz_rom_97[69] = 1'b0;
      zz_rom_97[70] = 1'b0;
      zz_rom_97[71] = 1'b0;
      zz_rom_97[72] = 1'b0;
      zz_rom_97[73] = 1'b0;
      zz_rom_97[74] = 1'b0;
      zz_rom_97[75] = 1'b0;
      zz_rom_97[76] = 1'b0;
      zz_rom_97[77] = 1'b0;
      zz_rom_97[78] = 1'b0;
      zz_rom_97[79] = 1'b0;
      zz_rom_97[80] = 1'b0;
      zz_rom_97[81] = 1'b0;
      zz_rom_97[82] = 1'b0;
      zz_rom_97[83] = 1'b0;
      zz_rom_97[84] = 1'b0;
      zz_rom_97[85] = 1'b0;
      zz_rom_97[86] = 1'b0;
      zz_rom_97[87] = 1'b0;
      zz_rom_97[88] = 1'b0;
      zz_rom_97[89] = 1'b0;
      zz_rom_97[90] = 1'b0;
      zz_rom_97[91] = 1'b0;
      zz_rom_97[92] = 1'b0;
      zz_rom_97[93] = 1'b0;
      zz_rom_97[94] = 1'b0;
      zz_rom_97[95] = 1'b0;
      zz_rom_97[96] = 1'b0;
      zz_rom_97[97] = 1'b0;
      zz_rom_97[98] = 1'b0;
      zz_rom_97[99] = 1'b0;
    end
  endfunction
  wire [99:0] _zz_98;
  function [99:0] zz_rom_98(input dummy);
    begin
      zz_rom_98[0] = 1'b0;
      zz_rom_98[1] = 1'b0;
      zz_rom_98[2] = 1'b0;
      zz_rom_98[3] = 1'b0;
      zz_rom_98[4] = 1'b0;
      zz_rom_98[5] = 1'b0;
      zz_rom_98[6] = 1'b0;
      zz_rom_98[7] = 1'b0;
      zz_rom_98[8] = 1'b0;
      zz_rom_98[9] = 1'b0;
      zz_rom_98[10] = 1'b0;
      zz_rom_98[11] = 1'b0;
      zz_rom_98[12] = 1'b0;
      zz_rom_98[13] = 1'b0;
      zz_rom_98[14] = 1'b0;
      zz_rom_98[15] = 1'b0;
      zz_rom_98[16] = 1'b0;
      zz_rom_98[17] = 1'b0;
      zz_rom_98[18] = 1'b0;
      zz_rom_98[19] = 1'b0;
      zz_rom_98[20] = 1'b0;
      zz_rom_98[21] = 1'b0;
      zz_rom_98[22] = 1'b0;
      zz_rom_98[23] = 1'b0;
      zz_rom_98[24] = 1'b0;
      zz_rom_98[25] = 1'b0;
      zz_rom_98[26] = 1'b0;
      zz_rom_98[27] = 1'b0;
      zz_rom_98[28] = 1'b0;
      zz_rom_98[29] = 1'b0;
      zz_rom_98[30] = 1'b0;
      zz_rom_98[31] = 1'b0;
      zz_rom_98[32] = 1'b0;
      zz_rom_98[33] = 1'b0;
      zz_rom_98[34] = 1'b0;
      zz_rom_98[35] = 1'b0;
      zz_rom_98[36] = 1'b1;
      zz_rom_98[37] = 1'b1;
      zz_rom_98[38] = 1'b1;
      zz_rom_98[39] = 1'b1;
      zz_rom_98[40] = 1'b1;
      zz_rom_98[41] = 1'b1;
      zz_rom_98[42] = 1'b1;
      zz_rom_98[43] = 1'b1;
      zz_rom_98[44] = 1'b1;
      zz_rom_98[45] = 1'b1;
      zz_rom_98[46] = 1'b1;
      zz_rom_98[47] = 1'b1;
      zz_rom_98[48] = 1'b1;
      zz_rom_98[49] = 1'b1;
      zz_rom_98[50] = 1'b1;
      zz_rom_98[51] = 1'b1;
      zz_rom_98[52] = 1'b1;
      zz_rom_98[53] = 1'b1;
      zz_rom_98[54] = 1'b1;
      zz_rom_98[55] = 1'b1;
      zz_rom_98[56] = 1'b1;
      zz_rom_98[57] = 1'b1;
      zz_rom_98[58] = 1'b1;
      zz_rom_98[59] = 1'b1;
      zz_rom_98[60] = 1'b1;
      zz_rom_98[61] = 1'b1;
      zz_rom_98[62] = 1'b1;
      zz_rom_98[63] = 1'b1;
      zz_rom_98[64] = 1'b1;
      zz_rom_98[65] = 1'b0;
      zz_rom_98[66] = 1'b0;
      zz_rom_98[67] = 1'b0;
      zz_rom_98[68] = 1'b0;
      zz_rom_98[69] = 1'b0;
      zz_rom_98[70] = 1'b0;
      zz_rom_98[71] = 1'b0;
      zz_rom_98[72] = 1'b0;
      zz_rom_98[73] = 1'b0;
      zz_rom_98[74] = 1'b0;
      zz_rom_98[75] = 1'b0;
      zz_rom_98[76] = 1'b0;
      zz_rom_98[77] = 1'b0;
      zz_rom_98[78] = 1'b0;
      zz_rom_98[79] = 1'b0;
      zz_rom_98[80] = 1'b0;
      zz_rom_98[81] = 1'b0;
      zz_rom_98[82] = 1'b0;
      zz_rom_98[83] = 1'b0;
      zz_rom_98[84] = 1'b0;
      zz_rom_98[85] = 1'b0;
      zz_rom_98[86] = 1'b0;
      zz_rom_98[87] = 1'b0;
      zz_rom_98[88] = 1'b0;
      zz_rom_98[89] = 1'b0;
      zz_rom_98[90] = 1'b0;
      zz_rom_98[91] = 1'b0;
      zz_rom_98[92] = 1'b0;
      zz_rom_98[93] = 1'b0;
      zz_rom_98[94] = 1'b0;
      zz_rom_98[95] = 1'b0;
      zz_rom_98[96] = 1'b0;
      zz_rom_98[97] = 1'b0;
      zz_rom_98[98] = 1'b0;
      zz_rom_98[99] = 1'b0;
    end
  endfunction
  wire [99:0] _zz_99;
  function [99:0] zz_rom_99(input dummy);
    begin
      zz_rom_99[0] = 1'b0;
      zz_rom_99[1] = 1'b0;
      zz_rom_99[2] = 1'b0;
      zz_rom_99[3] = 1'b0;
      zz_rom_99[4] = 1'b0;
      zz_rom_99[5] = 1'b0;
      zz_rom_99[6] = 1'b0;
      zz_rom_99[7] = 1'b0;
      zz_rom_99[8] = 1'b0;
      zz_rom_99[9] = 1'b0;
      zz_rom_99[10] = 1'b0;
      zz_rom_99[11] = 1'b0;
      zz_rom_99[12] = 1'b0;
      zz_rom_99[13] = 1'b0;
      zz_rom_99[14] = 1'b0;
      zz_rom_99[15] = 1'b0;
      zz_rom_99[16] = 1'b0;
      zz_rom_99[17] = 1'b0;
      zz_rom_99[18] = 1'b0;
      zz_rom_99[19] = 1'b0;
      zz_rom_99[20] = 1'b0;
      zz_rom_99[21] = 1'b0;
      zz_rom_99[22] = 1'b0;
      zz_rom_99[23] = 1'b0;
      zz_rom_99[24] = 1'b0;
      zz_rom_99[25] = 1'b0;
      zz_rom_99[26] = 1'b0;
      zz_rom_99[27] = 1'b0;
      zz_rom_99[28] = 1'b0;
      zz_rom_99[29] = 1'b0;
      zz_rom_99[30] = 1'b0;
      zz_rom_99[31] = 1'b0;
      zz_rom_99[32] = 1'b0;
      zz_rom_99[33] = 1'b0;
      zz_rom_99[34] = 1'b0;
      zz_rom_99[35] = 1'b0;
      zz_rom_99[36] = 1'b0;
      zz_rom_99[37] = 1'b0;
      zz_rom_99[38] = 1'b0;
      zz_rom_99[39] = 1'b0;
      zz_rom_99[40] = 1'b0;
      zz_rom_99[41] = 1'b1;
      zz_rom_99[42] = 1'b1;
      zz_rom_99[43] = 1'b1;
      zz_rom_99[44] = 1'b1;
      zz_rom_99[45] = 1'b1;
      zz_rom_99[46] = 1'b1;
      zz_rom_99[47] = 1'b1;
      zz_rom_99[48] = 1'b1;
      zz_rom_99[49] = 1'b1;
      zz_rom_99[50] = 1'b1;
      zz_rom_99[51] = 1'b1;
      zz_rom_99[52] = 1'b1;
      zz_rom_99[53] = 1'b1;
      zz_rom_99[54] = 1'b1;
      zz_rom_99[55] = 1'b1;
      zz_rom_99[56] = 1'b1;
      zz_rom_99[57] = 1'b1;
      zz_rom_99[58] = 1'b1;
      zz_rom_99[59] = 1'b1;
      zz_rom_99[60] = 1'b0;
      zz_rom_99[61] = 1'b0;
      zz_rom_99[62] = 1'b0;
      zz_rom_99[63] = 1'b0;
      zz_rom_99[64] = 1'b0;
      zz_rom_99[65] = 1'b0;
      zz_rom_99[66] = 1'b0;
      zz_rom_99[67] = 1'b0;
      zz_rom_99[68] = 1'b0;
      zz_rom_99[69] = 1'b0;
      zz_rom_99[70] = 1'b0;
      zz_rom_99[71] = 1'b0;
      zz_rom_99[72] = 1'b0;
      zz_rom_99[73] = 1'b0;
      zz_rom_99[74] = 1'b0;
      zz_rom_99[75] = 1'b0;
      zz_rom_99[76] = 1'b0;
      zz_rom_99[77] = 1'b0;
      zz_rom_99[78] = 1'b0;
      zz_rom_99[79] = 1'b0;
      zz_rom_99[80] = 1'b0;
      zz_rom_99[81] = 1'b0;
      zz_rom_99[82] = 1'b0;
      zz_rom_99[83] = 1'b0;
      zz_rom_99[84] = 1'b0;
      zz_rom_99[85] = 1'b0;
      zz_rom_99[86] = 1'b0;
      zz_rom_99[87] = 1'b0;
      zz_rom_99[88] = 1'b0;
      zz_rom_99[89] = 1'b0;
      zz_rom_99[90] = 1'b0;
      zz_rom_99[91] = 1'b0;
      zz_rom_99[92] = 1'b0;
      zz_rom_99[93] = 1'b0;
      zz_rom_99[94] = 1'b0;
      zz_rom_99[95] = 1'b0;
      zz_rom_99[96] = 1'b0;
      zz_rom_99[97] = 1'b0;
      zz_rom_99[98] = 1'b0;
      zz_rom_99[99] = 1'b0;
    end
  endfunction
  wire [99:0] _zz_100;

  assign _zz_x_offset = (io_x - x0);
  assign _zz_y_offset = (io_y - y0);
  assign _zz_when_shape_l120 = (x0 + diameter);
  assign _zz_when_shape_l120_1 = (y0 + diameter);
  always @(*) begin
    case(x_offset)
      7'b0000000 : _zz_xBits = rom_0;
      7'b0000001 : _zz_xBits = rom_1;
      7'b0000010 : _zz_xBits = rom_2;
      7'b0000011 : _zz_xBits = rom_3;
      7'b0000100 : _zz_xBits = rom_4;
      7'b0000101 : _zz_xBits = rom_5;
      7'b0000110 : _zz_xBits = rom_6;
      7'b0000111 : _zz_xBits = rom_7;
      7'b0001000 : _zz_xBits = rom_8;
      7'b0001001 : _zz_xBits = rom_9;
      7'b0001010 : _zz_xBits = rom_10;
      7'b0001011 : _zz_xBits = rom_11;
      7'b0001100 : _zz_xBits = rom_12;
      7'b0001101 : _zz_xBits = rom_13;
      7'b0001110 : _zz_xBits = rom_14;
      7'b0001111 : _zz_xBits = rom_15;
      7'b0010000 : _zz_xBits = rom_16;
      7'b0010001 : _zz_xBits = rom_17;
      7'b0010010 : _zz_xBits = rom_18;
      7'b0010011 : _zz_xBits = rom_19;
      7'b0010100 : _zz_xBits = rom_20;
      7'b0010101 : _zz_xBits = rom_21;
      7'b0010110 : _zz_xBits = rom_22;
      7'b0010111 : _zz_xBits = rom_23;
      7'b0011000 : _zz_xBits = rom_24;
      7'b0011001 : _zz_xBits = rom_25;
      7'b0011010 : _zz_xBits = rom_26;
      7'b0011011 : _zz_xBits = rom_27;
      7'b0011100 : _zz_xBits = rom_28;
      7'b0011101 : _zz_xBits = rom_29;
      7'b0011110 : _zz_xBits = rom_30;
      7'b0011111 : _zz_xBits = rom_31;
      7'b0100000 : _zz_xBits = rom_32;
      7'b0100001 : _zz_xBits = rom_33;
      7'b0100010 : _zz_xBits = rom_34;
      7'b0100011 : _zz_xBits = rom_35;
      7'b0100100 : _zz_xBits = rom_36;
      7'b0100101 : _zz_xBits = rom_37;
      7'b0100110 : _zz_xBits = rom_38;
      7'b0100111 : _zz_xBits = rom_39;
      7'b0101000 : _zz_xBits = rom_40;
      7'b0101001 : _zz_xBits = rom_41;
      7'b0101010 : _zz_xBits = rom_42;
      7'b0101011 : _zz_xBits = rom_43;
      7'b0101100 : _zz_xBits = rom_44;
      7'b0101101 : _zz_xBits = rom_45;
      7'b0101110 : _zz_xBits = rom_46;
      7'b0101111 : _zz_xBits = rom_47;
      7'b0110000 : _zz_xBits = rom_48;
      7'b0110001 : _zz_xBits = rom_49;
      7'b0110010 : _zz_xBits = rom_50;
      7'b0110011 : _zz_xBits = rom_51;
      7'b0110100 : _zz_xBits = rom_52;
      7'b0110101 : _zz_xBits = rom_53;
      7'b0110110 : _zz_xBits = rom_54;
      7'b0110111 : _zz_xBits = rom_55;
      7'b0111000 : _zz_xBits = rom_56;
      7'b0111001 : _zz_xBits = rom_57;
      7'b0111010 : _zz_xBits = rom_58;
      7'b0111011 : _zz_xBits = rom_59;
      7'b0111100 : _zz_xBits = rom_60;
      7'b0111101 : _zz_xBits = rom_61;
      7'b0111110 : _zz_xBits = rom_62;
      7'b0111111 : _zz_xBits = rom_63;
      7'b1000000 : _zz_xBits = rom_64;
      7'b1000001 : _zz_xBits = rom_65;
      7'b1000010 : _zz_xBits = rom_66;
      7'b1000011 : _zz_xBits = rom_67;
      7'b1000100 : _zz_xBits = rom_68;
      7'b1000101 : _zz_xBits = rom_69;
      7'b1000110 : _zz_xBits = rom_70;
      7'b1000111 : _zz_xBits = rom_71;
      7'b1001000 : _zz_xBits = rom_72;
      7'b1001001 : _zz_xBits = rom_73;
      7'b1001010 : _zz_xBits = rom_74;
      7'b1001011 : _zz_xBits = rom_75;
      7'b1001100 : _zz_xBits = rom_76;
      7'b1001101 : _zz_xBits = rom_77;
      7'b1001110 : _zz_xBits = rom_78;
      7'b1001111 : _zz_xBits = rom_79;
      7'b1010000 : _zz_xBits = rom_80;
      7'b1010001 : _zz_xBits = rom_81;
      7'b1010010 : _zz_xBits = rom_82;
      7'b1010011 : _zz_xBits = rom_83;
      7'b1010100 : _zz_xBits = rom_84;
      7'b1010101 : _zz_xBits = rom_85;
      7'b1010110 : _zz_xBits = rom_86;
      7'b1010111 : _zz_xBits = rom_87;
      7'b1011000 : _zz_xBits = rom_88;
      7'b1011001 : _zz_xBits = rom_89;
      7'b1011010 : _zz_xBits = rom_90;
      7'b1011011 : _zz_xBits = rom_91;
      7'b1011100 : _zz_xBits = rom_92;
      7'b1011101 : _zz_xBits = rom_93;
      7'b1011110 : _zz_xBits = rom_94;
      7'b1011111 : _zz_xBits = rom_95;
      7'b1100000 : _zz_xBits = rom_96;
      7'b1100001 : _zz_xBits = rom_97;
      7'b1100010 : _zz_xBits = rom_98;
      default : _zz_xBits = rom_99;
    endcase
  end

  assign x0 = 10'h0c8;
  assign y0 = 10'h12c;
  assign io_color_r = 4'b0000;
  assign io_color_g = 4'b0000;
  assign io_color_b = 4'b1111;
  assign diameter = 10'h064;
  assign _zz_1 = zz_rom_0(1'b0);
  always @(*) rom_0 = _zz_1;
  assign _zz_2 = zz_rom_1(1'b0);
  always @(*) rom_1 = _zz_2;
  assign _zz_3 = zz_rom_2(1'b0);
  always @(*) rom_2 = _zz_3;
  assign _zz_4 = zz_rom_3(1'b0);
  always @(*) rom_3 = _zz_4;
  assign _zz_5 = zz_rom_4(1'b0);
  always @(*) rom_4 = _zz_5;
  assign _zz_6 = zz_rom_5(1'b0);
  always @(*) rom_5 = _zz_6;
  assign _zz_7 = zz_rom_6(1'b0);
  always @(*) rom_6 = _zz_7;
  assign _zz_8 = zz_rom_7(1'b0);
  always @(*) rom_7 = _zz_8;
  assign _zz_9 = zz_rom_8(1'b0);
  always @(*) rom_8 = _zz_9;
  assign _zz_10 = zz_rom_9(1'b0);
  always @(*) rom_9 = _zz_10;
  assign _zz_11 = zz_rom_10(1'b0);
  always @(*) rom_10 = _zz_11;
  assign _zz_12 = zz_rom_11(1'b0);
  always @(*) rom_11 = _zz_12;
  assign _zz_13 = zz_rom_12(1'b0);
  always @(*) rom_12 = _zz_13;
  assign _zz_14 = zz_rom_13(1'b0);
  always @(*) rom_13 = _zz_14;
  assign _zz_15 = zz_rom_14(1'b0);
  always @(*) rom_14 = _zz_15;
  assign _zz_16 = zz_rom_15(1'b0);
  always @(*) rom_15 = _zz_16;
  assign _zz_17 = zz_rom_16(1'b0);
  always @(*) rom_16 = _zz_17;
  assign _zz_18 = zz_rom_17(1'b0);
  always @(*) rom_17 = _zz_18;
  assign _zz_19 = zz_rom_18(1'b0);
  always @(*) rom_18 = _zz_19;
  assign _zz_20 = zz_rom_19(1'b0);
  always @(*) rom_19 = _zz_20;
  assign _zz_21 = zz_rom_20(1'b0);
  always @(*) rom_20 = _zz_21;
  assign _zz_22 = zz_rom_21(1'b0);
  always @(*) rom_21 = _zz_22;
  assign _zz_23 = zz_rom_22(1'b0);
  always @(*) rom_22 = _zz_23;
  assign _zz_24 = zz_rom_23(1'b0);
  always @(*) rom_23 = _zz_24;
  assign _zz_25 = zz_rom_24(1'b0);
  always @(*) rom_24 = _zz_25;
  assign _zz_26 = zz_rom_25(1'b0);
  always @(*) rom_25 = _zz_26;
  assign _zz_27 = zz_rom_26(1'b0);
  always @(*) rom_26 = _zz_27;
  assign _zz_28 = zz_rom_27(1'b0);
  always @(*) rom_27 = _zz_28;
  assign _zz_29 = zz_rom_28(1'b0);
  always @(*) rom_28 = _zz_29;
  assign _zz_30 = zz_rom_29(1'b0);
  always @(*) rom_29 = _zz_30;
  assign _zz_31 = zz_rom_30(1'b0);
  always @(*) rom_30 = _zz_31;
  assign _zz_32 = zz_rom_31(1'b0);
  always @(*) rom_31 = _zz_32;
  assign _zz_33 = zz_rom_32(1'b0);
  always @(*) rom_32 = _zz_33;
  assign _zz_34 = zz_rom_33(1'b0);
  always @(*) rom_33 = _zz_34;
  assign _zz_35 = zz_rom_34(1'b0);
  always @(*) rom_34 = _zz_35;
  assign _zz_36 = zz_rom_35(1'b0);
  always @(*) rom_35 = _zz_36;
  assign _zz_37 = zz_rom_36(1'b0);
  always @(*) rom_36 = _zz_37;
  assign _zz_38 = zz_rom_37(1'b0);
  always @(*) rom_37 = _zz_38;
  assign _zz_39 = zz_rom_38(1'b0);
  always @(*) rom_38 = _zz_39;
  assign _zz_40 = zz_rom_39(1'b0);
  always @(*) rom_39 = _zz_40;
  assign _zz_41 = zz_rom_40(1'b0);
  always @(*) rom_40 = _zz_41;
  assign _zz_42 = zz_rom_41(1'b0);
  always @(*) rom_41 = _zz_42;
  assign _zz_43 = zz_rom_42(1'b0);
  always @(*) rom_42 = _zz_43;
  assign _zz_44 = zz_rom_43(1'b0);
  always @(*) rom_43 = _zz_44;
  assign _zz_45 = zz_rom_44(1'b0);
  always @(*) rom_44 = _zz_45;
  assign _zz_46 = zz_rom_45(1'b0);
  always @(*) rom_45 = _zz_46;
  assign _zz_47 = zz_rom_46(1'b0);
  always @(*) rom_46 = _zz_47;
  assign _zz_48 = zz_rom_47(1'b0);
  always @(*) rom_47 = _zz_48;
  assign _zz_49 = zz_rom_48(1'b0);
  always @(*) rom_48 = _zz_49;
  assign _zz_50 = zz_rom_49(1'b0);
  always @(*) rom_49 = _zz_50;
  assign _zz_51 = zz_rom_50(1'b0);
  always @(*) rom_50 = _zz_51;
  assign _zz_52 = zz_rom_51(1'b0);
  always @(*) rom_51 = _zz_52;
  assign _zz_53 = zz_rom_52(1'b0);
  always @(*) rom_52 = _zz_53;
  assign _zz_54 = zz_rom_53(1'b0);
  always @(*) rom_53 = _zz_54;
  assign _zz_55 = zz_rom_54(1'b0);
  always @(*) rom_54 = _zz_55;
  assign _zz_56 = zz_rom_55(1'b0);
  always @(*) rom_55 = _zz_56;
  assign _zz_57 = zz_rom_56(1'b0);
  always @(*) rom_56 = _zz_57;
  assign _zz_58 = zz_rom_57(1'b0);
  always @(*) rom_57 = _zz_58;
  assign _zz_59 = zz_rom_58(1'b0);
  always @(*) rom_58 = _zz_59;
  assign _zz_60 = zz_rom_59(1'b0);
  always @(*) rom_59 = _zz_60;
  assign _zz_61 = zz_rom_60(1'b0);
  always @(*) rom_60 = _zz_61;
  assign _zz_62 = zz_rom_61(1'b0);
  always @(*) rom_61 = _zz_62;
  assign _zz_63 = zz_rom_62(1'b0);
  always @(*) rom_62 = _zz_63;
  assign _zz_64 = zz_rom_63(1'b0);
  always @(*) rom_63 = _zz_64;
  assign _zz_65 = zz_rom_64(1'b0);
  always @(*) rom_64 = _zz_65;
  assign _zz_66 = zz_rom_65(1'b0);
  always @(*) rom_65 = _zz_66;
  assign _zz_67 = zz_rom_66(1'b0);
  always @(*) rom_66 = _zz_67;
  assign _zz_68 = zz_rom_67(1'b0);
  always @(*) rom_67 = _zz_68;
  assign _zz_69 = zz_rom_68(1'b0);
  always @(*) rom_68 = _zz_69;
  assign _zz_70 = zz_rom_69(1'b0);
  always @(*) rom_69 = _zz_70;
  assign _zz_71 = zz_rom_70(1'b0);
  always @(*) rom_70 = _zz_71;
  assign _zz_72 = zz_rom_71(1'b0);
  always @(*) rom_71 = _zz_72;
  assign _zz_73 = zz_rom_72(1'b0);
  always @(*) rom_72 = _zz_73;
  assign _zz_74 = zz_rom_73(1'b0);
  always @(*) rom_73 = _zz_74;
  assign _zz_75 = zz_rom_74(1'b0);
  always @(*) rom_74 = _zz_75;
  assign _zz_76 = zz_rom_75(1'b0);
  always @(*) rom_75 = _zz_76;
  assign _zz_77 = zz_rom_76(1'b0);
  always @(*) rom_76 = _zz_77;
  assign _zz_78 = zz_rom_77(1'b0);
  always @(*) rom_77 = _zz_78;
  assign _zz_79 = zz_rom_78(1'b0);
  always @(*) rom_78 = _zz_79;
  assign _zz_80 = zz_rom_79(1'b0);
  always @(*) rom_79 = _zz_80;
  assign _zz_81 = zz_rom_80(1'b0);
  always @(*) rom_80 = _zz_81;
  assign _zz_82 = zz_rom_81(1'b0);
  always @(*) rom_81 = _zz_82;
  assign _zz_83 = zz_rom_82(1'b0);
  always @(*) rom_82 = _zz_83;
  assign _zz_84 = zz_rom_83(1'b0);
  always @(*) rom_83 = _zz_84;
  assign _zz_85 = zz_rom_84(1'b0);
  always @(*) rom_84 = _zz_85;
  assign _zz_86 = zz_rom_85(1'b0);
  always @(*) rom_85 = _zz_86;
  assign _zz_87 = zz_rom_86(1'b0);
  always @(*) rom_86 = _zz_87;
  assign _zz_88 = zz_rom_87(1'b0);
  always @(*) rom_87 = _zz_88;
  assign _zz_89 = zz_rom_88(1'b0);
  always @(*) rom_88 = _zz_89;
  assign _zz_90 = zz_rom_89(1'b0);
  always @(*) rom_89 = _zz_90;
  assign _zz_91 = zz_rom_90(1'b0);
  always @(*) rom_90 = _zz_91;
  assign _zz_92 = zz_rom_91(1'b0);
  always @(*) rom_91 = _zz_92;
  assign _zz_93 = zz_rom_92(1'b0);
  always @(*) rom_92 = _zz_93;
  assign _zz_94 = zz_rom_93(1'b0);
  always @(*) rom_93 = _zz_94;
  assign _zz_95 = zz_rom_94(1'b0);
  always @(*) rom_94 = _zz_95;
  assign _zz_96 = zz_rom_95(1'b0);
  always @(*) rom_95 = _zz_96;
  assign _zz_97 = zz_rom_96(1'b0);
  always @(*) rom_96 = _zz_97;
  assign _zz_98 = zz_rom_97(1'b0);
  always @(*) rom_97 = _zz_98;
  assign _zz_99 = zz_rom_98(1'b0);
  always @(*) rom_98 = _zz_99;
  assign _zz_100 = zz_rom_99(1'b0);
  always @(*) rom_99 = _zz_100;
  assign x_offset = _zz_x_offset[6:0];
  assign y_offset = _zz_y_offset[6:0];
  assign xBits = _zz_xBits;
  assign when_shape_l120 = ((((x0 <= io_x) && (io_x < _zz_when_shape_l120)) && (y0 <= io_y)) && (io_y < _zz_when_shape_l120_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      io_inside <= 1'b0;
    end else begin
      if(when_shape_l120) begin
        io_inside <= xBits[y_offset];
      end else begin
        io_inside <= 1'b0;
      end
    end
  end


endmodule

module square (
  input      [9:0]    io_x,
  input      [9:0]    io_y,
  output reg          io_inside,
  output     [3:0]    io_color_r,
  output     [3:0]    io_color_g,
  output     [3:0]    io_color_b,
  input               clk,
  input               reset
);

  wire       [9:0]    _zz_when_shape_l88;
  wire       [9:0]    _zz_when_shape_l88_1;
  wire       [9:0]    x0;
  wire       [9:0]    y0;
  wire       [9:0]    x_width;
  wire       [9:0]    y_height;
  wire                when_shape_l88;

  assign _zz_when_shape_l88 = (x0 + x_width);
  assign _zz_when_shape_l88_1 = (y0 + y_height);
  assign x0 = 10'h06e;
  assign y0 = 10'h014;
  assign io_color_r = 4'b0000;
  assign io_color_g = 4'b1111;
  assign io_color_b = 4'b0000;
  assign x_width = 10'h03c;
  assign y_height = 10'h03c;
  assign when_shape_l88 = ((((x0 <= io_x) && (io_x < _zz_when_shape_l88)) && (y0 <= io_y)) && (io_y < _zz_when_shape_l88_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      io_inside <= 1'b0;
    end else begin
      if(when_shape_l88) begin
        io_inside <= 1'b1;
      end else begin
        io_inside <= 1'b0;
      end
    end
  end


endmodule

module rectangle (
  input      [9:0]    io_x,
  input      [9:0]    io_y,
  output reg          io_inside,
  output     [3:0]    io_color_r,
  output     [3:0]    io_color_g,
  output     [3:0]    io_color_b,
  input               clk,
  input               reset
);

  wire       [9:0]    _zz_when_shape_l88;
  wire       [9:0]    _zz_when_shape_l88_1;
  wire       [9:0]    x0;
  wire       [9:0]    y0;
  wire       [9:0]    x_width;
  wire       [9:0]    y_height;
  wire                when_shape_l88;

  assign _zz_when_shape_l88 = (x0 + x_width);
  assign _zz_when_shape_l88_1 = (y0 + y_height);
  assign x0 = 10'h00a;
  assign y0 = 10'h014;
  assign io_color_r = 4'b1111;
  assign io_color_g = 4'b0000;
  assign io_color_b = 4'b0000;
  assign x_width = 10'h014;
  assign y_height = 10'h078;
  assign when_shape_l88 = ((((x0 <= io_x) && (io_x < _zz_when_shape_l88)) && (y0 <= io_y)) && (io_y < _zz_when_shape_l88_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      io_inside <= 1'b0;
    end else begin
      if(when_shape_l88) begin
        io_inside <= 1'b1;
      end else begin
        io_inside <= 1'b0;
      end
    end
  end


endmodule
